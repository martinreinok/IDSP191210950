
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_MAP1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type SIGNED is array (INTEGER range <>) of std_logic;

end CONV_PACK_MAP1;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_MAP1.all;

architecture flat_rtl_none_10 of MAP1 is

   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4M1D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal arx_i1_reg_7_port, arx_i1_reg_6_port, arx_i1_reg_5_port, 
      arx_i1_reg_4_port, arx_i1_reg_3_port, arx_i1_reg_2_port, 
      arx_i1_reg_1_port, arx_i1_reg_0_port, arx_r1_reg_14_port, 
      arx_r1_reg_13_port, arx_r1_reg_12_port, arx_r1_reg_11_port, 
      arx_r1_reg_10_port, arx_r1_reg_9_port, arx_r1_reg_8_port, 
      arx_r1_reg_7_port, arx_r1_reg_6_port, arx_r1_reg_5_port, 
      arx_r1_reg_4_port, arx_r1_reg_3_port, arx_r1_reg_2_port, 
      arx_r1_reg_1_port, arx_r1_reg_0_port, arx_r2_reg_14_port, 
      arx_r2_reg_13_port, arx_r2_reg_12_port, arx_r2_reg_11_port, 
      arx_r2_reg_10_port, arx_r2_reg_9_port, arx_r2_reg_8_port, 
      arx_r2_reg_7_port, arx_r2_reg_6_port, arx_r2_reg_5_port, 
      arx_r2_reg_4_port, arx_r2_reg_3_port, arx_r2_reg_2_port, 
      arx_r2_reg_1_port, arx_r2_reg_0_port, arx_state_reg_2_port, 
      arx_state_reg_1_port, arx_state_reg_0_port, m_in_l_4, m_in_l_0, 
      m_in_r_7_port, m_in_r_6_port, m_in_r_5_port, m_in_r_4_port, m_in_r_3_port
      , m_in_r_2_port, m_in_r_1_port, m_in_r_0_port, m_out_14_port, 
      m_out_13_port, m_out_12_port, m_out_11_port, m_out_10_port, m_out_9_port,
      m_out_8_port, m_out_7_port, m_out_6_port, m_out_5_port, m_out_4_port, 
      m_out_3_port, m_out_2_port, m_out_1_port, m_out_0_port, m2_in_l_5_port, 
      m2_in_l_3_port, m2_in_r_7_port, m2_in_r_6_port, m2_in_r_5_port, 
      m2_in_r_4_port, m2_in_r_3_port, m2_in_r_2_port, m2_in_r_1_port, 
      m2_in_r_0_port, m2_out_14_port, m2_out_13_port, m2_out_12_port, 
      m2_out_11_port, m2_out_10_port, m2_out_9_port, m2_out_8_port, 
      m2_out_7_port, m2_out_6_port, m2_out_5_port, m2_out_4_port, m2_out_3_port
      , m2_out_2_port, m2_out_1_port, m2_out_0_port, a_in_l_14_port, 
      a_in_l_13_port, a_in_l_12_port, a_in_l_11_port, a_in_l_10_port, 
      a_in_l_9_port, a_in_l_8_port, a_in_l_7_port, a_in_l_6_port, a_in_l_5_port
      , a_in_l_4_port, a_in_l_3_port, a_in_l_2_port, a_in_l_1_port, 
      a_in_l_0_port, a_in_r_14_port, a_in_r_13_port, a_in_r_12_port, 
      a_in_r_11_port, a_in_r_10_port, a_in_r_9_port, a_in_r_8_port, 
      a_in_r_7_port, a_in_r_6_port, a_in_r_5_port, a_in_r_4_port, a_in_r_3_port
      , a_in_r_2_port, a_in_r_1_port, a_in_r_0_port, a_out_7_port, a_out_6_port
      , a_out_5_port, a_out_4_port, a_out_3_port, a_out_2_port, a_out_1_port, 
      a_out_0_port, state_2_port, state_1_port, state_0_port, N44, N45, N46, 
      N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N144, 
      N145, N146, N147, N148, N149, N150, N151, N152, net1366, n62, n63, n64, 
      n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n104, n105, n106, n107, n108, 
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, add_416_C204_rn_carry_1_port, add_416_C204_rn_carry_2_port, 
      add_416_C204_rn_carry_3_port, add_416_C204_rn_carry_4_port, 
      add_416_C204_rn_carry_5_port, add_416_C204_rn_carry_6_port, 
      add_416_C204_rn_carry_7_port, n175, n176, n177, n178, n179, n180, n181, 
      n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
      n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, 
      n206, n207, n208, n209, n210, n211, n212, n_1012, n_1013, n_1014, n_1015,
      n_1016, n_1017, n_1018, n_1019, n_1020, add_204_n9, add_204_n8, 
      add_204_n7, add_204_n6, add_204_n5, add_204_n4, add_204_n3, add_204_n2, 
      add_204_n1, add_204_carry_6_port, add_204_carry_7_port, 
      add_204_carry_8_port, add_204_carry_9_port, add_204_carry_10_port, 
      add_204_carry_11_port, add_204_carry_12_port, add_204_carry_13_port, 
      add_204_carry_14_port, mult_203_n241, mult_203_n240, mult_203_n239, 
      mult_203_n238, mult_203_n237, mult_203_n236, mult_203_n235, mult_203_n234
      , mult_203_n233, mult_203_n232, mult_203_n231, mult_203_n230, 
      mult_203_n229, mult_203_n228, mult_203_n227, mult_203_n226, mult_203_n225
      , mult_203_n224, mult_203_n223, mult_203_n222, mult_203_n221, 
      mult_203_n220, mult_203_n219, mult_203_n218, mult_203_n217, mult_203_n216
      , mult_203_n215, mult_203_n214, mult_203_n213, mult_203_n212, 
      mult_203_n211, mult_203_n210, mult_203_n209, mult_203_n208, mult_203_n207
      , mult_203_n206, mult_203_n205, mult_203_n204, mult_203_n203, 
      mult_203_n202, mult_203_n201, mult_203_n200, mult_203_n199, mult_203_n198
      , mult_203_n197, mult_203_n196, mult_203_n195, mult_203_n194, 
      mult_203_n92, mult_203_n91, mult_203_n90, mult_203_n89, mult_203_n88, 
      mult_203_n87, mult_203_n86, mult_203_n85, mult_203_n83, mult_203_n82, 
      mult_203_n81, mult_203_n80, mult_203_n79, mult_203_n77, mult_203_n76, 
      mult_203_n75, mult_203_n74, mult_203_n73, mult_203_n72, mult_203_n71, 
      mult_203_n70, mult_203_n69, mult_203_n68, mult_203_n67, mult_203_n65, 
      mult_203_n64, mult_203_n63, mult_203_n62, mult_203_n60, mult_203_n59, 
      mult_203_n58, mult_203_n57, mult_203_n56, mult_203_n55, mult_203_n54, 
      mult_203_n53, mult_203_n52, mult_203_n51, mult_203_n50, mult_203_n49, 
      mult_203_n48, mult_203_n47, mult_203_n46, mult_203_n45, mult_203_n44, 
      mult_203_n43, mult_203_n42, mult_203_n41, mult_203_n40, mult_203_n39, 
      mult_203_n38, mult_203_n37, mult_203_n36, mult_203_n35, mult_203_n34, 
      mult_203_n33, mult_203_n31, mult_203_n30, mult_203_n29, mult_203_n28, 
      mult_203_n27, mult_203_n26, mult_203_n25, mult_203_n24, mult_203_n23, 
      mult_203_n21, mult_203_n20, mult_203_n19, mult_203_n18, mult_203_n17, 
      mult_203_n16, mult_203_n14, mult_203_n12, mult_203_n11, mult_203_n10, 
      mult_203_n9, mult_203_n8, mult_203_n7, mult_203_n6, mult_203_n5, 
      mult_203_n4, mult_203_n3, mult_203_n2, mult_202_n181, mult_202_n180, 
      mult_202_n179, mult_202_n178, mult_202_n177, mult_202_n176, mult_202_n175
      , mult_202_n174, mult_202_n173, mult_202_n172, mult_202_n171, 
      mult_202_n170, mult_202_n169, mult_202_n168, mult_202_n167, mult_202_n115
      , mult_202_n114, mult_202_n113, mult_202_n112, mult_202_n111, 
      mult_202_n110, mult_202_n109, mult_202_n108, mult_202_n107, mult_202_n106
      , mult_202_n105, mult_202_n104, mult_202_n103, mult_202_n102, 
      mult_202_n101, mult_202_n100, mult_202_n99, mult_202_n98, mult_202_n97, 
      mult_202_n96, mult_202_n94, mult_202_n93, mult_202_n92, mult_202_n91, 
      mult_202_n90, mult_202_n89, mult_202_n88, mult_202_n87, mult_202_n86, 
      mult_202_n85, mult_202_n84, mult_202_n82, mult_202_n81, mult_202_n80, 
      mult_202_n79, mult_202_n78, mult_202_n77, mult_202_n76, mult_202_n75, 
      mult_202_n74, mult_202_n73, mult_202_n72, mult_202_n70, mult_202_n69, 
      mult_202_n68, mult_202_n67, mult_202_n66, mult_202_n65, mult_202_n64, 
      mult_202_n63, mult_202_n62, mult_202_n61, mult_202_n60, mult_202_n59, 
      mult_202_n58, mult_202_n57, mult_202_n56, mult_202_n55, mult_202_n54, 
      mult_202_n53, mult_202_n52, mult_202_n51, mult_202_n50, mult_202_n49, 
      mult_202_n48, mult_202_n47, mult_202_n46, mult_202_n45, mult_202_n44, 
      mult_202_n43, mult_202_n42, mult_202_n41, mult_202_n40, mult_202_n39, 
      mult_202_n38, mult_202_n36, mult_202_n35, mult_202_n34, mult_202_n33, 
      mult_202_n32, mult_202_n31, mult_202_n30, mult_202_n29, mult_202_n28, 
      mult_202_n27, mult_202_n26, mult_202_n25, mult_202_n24, mult_202_n23, 
      mult_202_n22, mult_202_n21, mult_202_n20, mult_202_n18, mult_202_n17, 
      mult_202_n16, mult_202_n15, mult_202_n14, mult_202_n13, mult_202_n12, 
      mult_202_n11, mult_202_n10, mult_202_n9, mult_202_n8, mult_202_n7, 
      mult_202_n6, mult_202_n5, mult_202_n4, mult_202_n3, mult_202_n2 : 
      std_logic;

begin
   
   U103 : OAI21D1 port map( A1 => n65, A2 => n212, B => n66, Z => n104);
   U104 : AOI22D1 port map( A1 => a_out_7_port, A2 => n67, B1 => m2_out_14_port
                           , B2 => n68, Z => n66);
   U105 : OAI21D1 port map( A1 => n65, A2 => n211, B => n69, Z => n105);
   U106 : AOI22D1 port map( A1 => a_out_6_port, A2 => n67, B1 => m2_out_13_port
                           , B2 => n68, Z => n69);
   U107 : OAI21D1 port map( A1 => n65, A2 => n210, B => n70, Z => n106);
   U108 : AOI22D1 port map( A1 => a_out_5_port, A2 => n67, B1 => m2_out_12_port
                           , B2 => n68, Z => n70);
   U109 : OAI21D1 port map( A1 => n65, A2 => n209, B => n71, Z => n107);
   U110 : AOI22D1 port map( A1 => a_out_4_port, A2 => n67, B1 => m2_out_11_port
                           , B2 => n68, Z => n71);
   U111 : OAI21D1 port map( A1 => n65, A2 => n208, B => n72, Z => n108);
   U112 : AOI22D1 port map( A1 => a_out_3_port, A2 => n67, B1 => m2_out_10_port
                           , B2 => n68, Z => n72);
   U113 : OAI21D1 port map( A1 => n65, A2 => n207, B => n73, Z => n109);
   U114 : AOI22D1 port map( A1 => a_out_2_port, A2 => n67, B1 => m2_out_9_port,
                           B2 => n68, Z => n73);
   U115 : OAI21D1 port map( A1 => n65, A2 => n206, B => n74, Z => n110);
   U116 : AOI22D1 port map( A1 => a_out_1_port, A2 => n67, B1 => m2_out_8_port,
                           B2 => n68, Z => n74);
   U117 : OAI21D1 port map( A1 => n65, A2 => n205, B => n75, Z => n111);
   U118 : AOI22D1 port map( A1 => a_out_0_port, A2 => n67, B1 => m2_out_7_port,
                           B2 => n68, Z => n75);
   U119 : OAI22M10D1 port map( A1 => m2_out_6_port, A2 => n176, B1 => n65, B2 
                           => n198, Z => n112);
   U120 : OAI22M10D1 port map( A1 => m2_out_5_port, A2 => n176, B1 => n65, B2 
                           => n199, Z => n113);
   U121 : OAI22M10D1 port map( A1 => m2_out_4_port, A2 => n176, B1 => n65, B2 
                           => n200, Z => n114);
   U122 : OAI22M10D1 port map( A1 => m2_out_3_port, A2 => n176, B1 => n65, B2 
                           => n201, Z => n115);
   U123 : OAI22M10D1 port map( A1 => m2_out_2_port, A2 => n176, B1 => n65, B2 
                           => n202, Z => n116);
   U124 : OAI22M10D1 port map( A1 => m2_out_1_port, A2 => n176, B1 => n65, B2 
                           => n203, Z => n117);
   U125 : OAI22M10D1 port map( A1 => m2_out_0_port, A2 => n176, B1 => n65, B2 
                           => n204, Z => n118);
   U126 : OAI21D1 port map( A1 => n80, A2 => n197, B => n81, Z => n119);
   U127 : AOI22D1 port map( A1 => m_out_0_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_0_port, Z => n81);
   U128 : OAI21D1 port map( A1 => n80, A2 => n196, B => n82, Z => n120);
   U129 : AOI22D1 port map( A1 => m_out_1_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_1_port, Z => n82);
   U130 : OAI21D1 port map( A1 => n80, A2 => n195, B => n83, Z => n121);
   U131 : AOI22D1 port map( A1 => m_out_2_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_2_port, Z => n83);
   U132 : OAI21D1 port map( A1 => n80, A2 => n194, B => n84, Z => n122);
   U133 : AOI22D1 port map( A1 => m_out_3_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_3_port, Z => n84);
   U134 : OAI21D1 port map( A1 => n80, A2 => n193, B => n85, Z => n123);
   U135 : AOI22D1 port map( A1 => m_out_4_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_4_port, Z => n85);
   U136 : OAI21D1 port map( A1 => n80, A2 => n192, B => n86, Z => n124);
   U137 : AOI22D1 port map( A1 => m_out_5_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_5_port, Z => n86);
   U138 : OAI21D1 port map( A1 => n80, A2 => n191, B => n87, Z => n125);
   U139 : AOI22D1 port map( A1 => m_out_6_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_6_port, Z => n87);
   U140 : OAI21D1 port map( A1 => n80, A2 => n190, B => n88, Z => n126);
   U141 : AOI22D1 port map( A1 => m_out_7_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_7_port, Z => n88);
   U142 : OAI21D1 port map( A1 => n80, A2 => n189, B => n89, Z => n127);
   U143 : AOI22D1 port map( A1 => m_out_8_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_8_port, Z => n89);
   U144 : OAI21D1 port map( A1 => n80, A2 => n188, B => n90, Z => n128);
   U145 : AOI22D1 port map( A1 => m_out_9_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_9_port, Z => n90);
   U146 : OAI21D1 port map( A1 => n80, A2 => n187, B => n91, Z => n129);
   U147 : AOI22D1 port map( A1 => m_out_10_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_10_port, Z => n91);
   U148 : OAI21D1 port map( A1 => n80, A2 => n186, B => n92, Z => n130);
   U149 : AOI22D1 port map( A1 => m_out_11_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_11_port, Z => n92);
   U150 : OAI21D1 port map( A1 => n80, A2 => n185, B => n93, Z => n131);
   U151 : AOI22D1 port map( A1 => m_out_12_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_12_port, Z => n93);
   U152 : OAI21D1 port map( A1 => n80, A2 => n184, B => n94, Z => n132);
   U153 : AOI22D1 port map( A1 => m_out_13_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_13_port, Z => n94);
   U154 : OAI21D1 port map( A1 => n80, A2 => n183, B => n95, Z => n133);
   U155 : AOI22D1 port map( A1 => m_out_14_port, A2 => n68, B1 => n77, B2 => 
                           m2_out_14_port, Z => n95);
   U156 : OAI22M10D1 port map( A1 => arx_i1_reg_2_port, A2 => n96, B1 => n102, 
                           B2 => n188, Z => a_in_l_9_port);
   U157 : OAI22M10D1 port map( A1 => arx_i1_reg_1_port, A2 => n96, B1 => n102, 
                           B2 => n189, Z => a_in_l_8_port);
   U158 : OAI22M10D1 port map( A1 => arx_i1_reg_0_port, A2 => n96, B1 => n102, 
                           B2 => n190, Z => a_in_l_7_port);
   U159 : OAI22M10D1 port map( A1 => arx_i1_reg_7_port, A2 => n96, B1 => n102, 
                           B2 => n183, Z => a_in_l_14_port);
   U160 : OAI22M10D1 port map( A1 => arx_i1_reg_6_port, A2 => n96, B1 => n102, 
                           B2 => n184, Z => a_in_l_13_port);
   U161 : OAI22M10D1 port map( A1 => arx_i1_reg_5_port, A2 => n96, B1 => n102, 
                           B2 => n185, Z => a_in_l_12_port);
   U162 : OAI22M10D1 port map( A1 => arx_i1_reg_4_port, A2 => n96, B1 => n102, 
                           B2 => n186, Z => a_in_l_11_port);
   U163 : OAI22M10D1 port map( A1 => arx_i1_reg_3_port, A2 => n96, B1 => n102, 
                           B2 => n187, Z => a_in_l_10_port);
   arx_r2_reg_reg_14 : DFFRPQ1 port map( D => n104, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_14_port);
   arx_r1_reg_reg_14 : DFFRPQ1 port map( D => n133, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_14_port);
   arx_i1_reg_reg_7 : DFERPQ1 port map( D => data_in(7), CEB => n97, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_7_port);
   arx_r2_reg_reg_13 : DFFRPQ1 port map( D => n105, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_13_port);
   arx_r1_reg_reg_13 : DFFRPQ1 port map( D => n132, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_13_port);
   arx_i1_reg_reg_6 : DFERPQ1 port map( D => data_in(6), CEB => n97, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_6_port);
   arx_r2_reg_reg_12 : DFFRPQ1 port map( D => n106, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_12_port);
   arx_r1_reg_reg_12 : DFFRPQ1 port map( D => n131, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_12_port);
   arx_i1_reg_reg_5 : DFERPQ1 port map( D => data_in(5), CEB => n97, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_5_port);
   arx_r2_reg_reg_11 : DFFRPQ1 port map( D => n107, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_11_port);
   arx_r1_reg_reg_11 : DFFRPQ1 port map( D => n130, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_11_port);
   arx_i1_reg_reg_4 : DFERPQ1 port map( D => data_in(4), CEB => n97, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_4_port);
   arx_r2_reg_reg_10 : DFFRPQ1 port map( D => n108, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_10_port);
   arx_r1_reg_reg_10 : DFFRPQ1 port map( D => n129, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_10_port);
   arx_i1_reg_reg_3 : DFERPQ1 port map( D => data_in(3), CEB => n97, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_3_port);
   arx_r2_reg_reg_9 : DFFRPQ1 port map( D => n109, CK => clock, RB => resetn, Q
                           => arx_r2_reg_9_port);
   arx_r1_reg_reg_9 : DFFRPQ1 port map( D => n128, CK => clock, RB => resetn, Q
                           => arx_r1_reg_9_port);
   arx_i1_reg_reg_2 : DFERPQ1 port map( D => data_in(2), CEB => n97, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_2_port);
   arx_r2_reg_reg_8 : DFFRPQ1 port map( D => n110, CK => clock, RB => resetn, Q
                           => arx_r2_reg_8_port);
   arx_r1_reg_reg_8 : DFFRPQ1 port map( D => n127, CK => clock, RB => resetn, Q
                           => arx_r1_reg_8_port);
   arx_i1_reg_reg_1 : DFERPQ1 port map( D => data_in(1), CEB => n97, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_1_port);
   arx_r2_reg_reg_7 : DFFRPQ1 port map( D => n111, CK => clock, RB => resetn, Q
                           => arx_r2_reg_7_port);
   arx_r1_reg_reg_7 : DFFRPQ1 port map( D => n126, CK => clock, RB => resetn, Q
                           => arx_r1_reg_7_port);
   arx_i1_reg_reg_0 : DFERPQ1 port map( D => data_in(0), CEB => n97, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_0_port);
   arx_r1_reg_reg_6 : DFFRPQ1 port map( D => n125, CK => clock, RB => resetn, Q
                           => arx_r1_reg_6_port);
   arx_r2_reg_reg_6 : DFFRPQ1 port map( D => n112, CK => clock, RB => resetn, Q
                           => arx_r2_reg_6_port);
   arx_r2_reg_reg_5 : DFFRPQ1 port map( D => n113, CK => clock, RB => resetn, Q
                           => arx_r2_reg_5_port);
   arx_r1_reg_reg_5 : DFFRPQ1 port map( D => n124, CK => clock, RB => resetn, Q
                           => arx_r1_reg_5_port);
   arx_r2_reg_reg_4 : DFFRPQ1 port map( D => n114, CK => clock, RB => resetn, Q
                           => arx_r2_reg_4_port);
   arx_r1_reg_reg_4 : DFFRPQ1 port map( D => n123, CK => clock, RB => resetn, Q
                           => arx_r1_reg_4_port);
   arx_r2_reg_reg_3 : DFFRPQ1 port map( D => n115, CK => clock, RB => resetn, Q
                           => arx_r2_reg_3_port);
   arx_r1_reg_reg_3 : DFFRPQ1 port map( D => n122, CK => clock, RB => resetn, Q
                           => arx_r1_reg_3_port);
   arx_d1_reg_reg_14 : DFERPQ1 port map( D => a_out_7_port, CEB => n64, CK => 
                           clock, RB => resetn, Q => N51);
   arx_r2_reg_reg_2 : DFFRPQ1 port map( D => n116, CK => clock, RB => resetn, Q
                           => arx_r2_reg_2_port);
   arx_r1_reg_reg_2 : DFFRPQ1 port map( D => n121, CK => clock, RB => resetn, Q
                           => arx_r1_reg_2_port);
   arx_d2_reg_reg_14 : DFERPQ1 port map( D => N51, CEB => n64, CK => clock, RB 
                           => resetn, Q => N59);
   arx_r2_reg_reg_0 : DFFRPQ1 port map( D => n118, CK => clock, RB => resetn, Q
                           => arx_r2_reg_0_port);
   arx_r1_reg_reg_0 : DFFRPQ1 port map( D => n119, CK => clock, RB => resetn, Q
                           => arx_r1_reg_0_port);
   arx_d1_reg_reg_13 : DFERPQ1 port map( D => a_out_6_port, CEB => n64, CK => 
                           clock, RB => resetn, Q => N50);
   arx_r1_reg_reg_1 : DFFRPQ1 port map( D => n120, CK => clock, RB => resetn, Q
                           => arx_r1_reg_1_port);
   arx_r2_reg_reg_1 : DFFRPQ1 port map( D => n117, CK => clock, RB => resetn, Q
                           => arx_r2_reg_1_port);
   arx_d1_reg_reg_12 : DFERPQ1 port map( D => a_out_5_port, CEB => n64, CK => 
                           clock, RB => resetn, Q => N49);
   arx_d2_reg_reg_13 : DFERPQ1 port map( D => N50, CEB => n64, CK => clock, RB 
                           => resetn, Q => N58);
   arx_d1_reg_reg_11 : DFERPQ1 port map( D => a_out_4_port, CEB => n64, CK => 
                           clock, RB => resetn, Q => N48);
   arx_d2_reg_reg_12 : DFERPQ1 port map( D => N49, CEB => n64, CK => clock, RB 
                           => resetn, Q => N57);
   arx_d1_reg_reg_9 : DFERPQ1 port map( D => a_out_2_port, CEB => n64, CK => 
                           clock, RB => resetn, Q => N46);
   arx_d1_reg_reg_8 : DFERPQ1 port map( D => a_out_1_port, CEB => n64, CK => 
                           clock, RB => resetn, Q => N45);
   arx_d1_reg_reg_10 : DFERPQ1 port map( D => a_out_3_port, CEB => n64, CK => 
                           clock, RB => resetn, Q => N47);
   arx_d1_reg_reg_7 : DFERPQ1 port map( D => a_out_0_port, CEB => n64, CK => 
                           clock, RB => resetn, Q => N44);
   arx_d2_reg_reg_11 : DFERPQ1 port map( D => N48, CEB => n64, CK => clock, RB 
                           => resetn, Q => N56);
   arx_d2_reg_reg_9 : DFERPQ1 port map( D => N46, CEB => n64, CK => clock, RB 
                           => resetn, Q => N54);
   arx_d2_reg_reg_8 : DFERPQ1 port map( D => N45, CEB => n64, CK => clock, RB 
                           => resetn, Q => N53);
   arx_d2_reg_reg_10 : DFERPQ1 port map( D => N47, CEB => n64, CK => clock, RB 
                           => resetn, Q => N55);
   arx_d2_reg_reg_7 : DFERPQ1 port map( D => N44, CEB => n64, CK => clock, RB 
                           => resetn, Q => N52);
   arx_state_reg_reg_0 : DFFRPQ1 port map( D => state_0_port, CK => clock, RB 
                           => resetn, Q => arx_state_reg_0_port);
   arx_state_reg_reg_1 : DFFRPQ1 port map( D => state_1_port, CK => clock, RB 
                           => resetn, Q => arx_state_reg_1_port);
   arx_state_reg_reg_2 : DFFRPQ1 port map( D => state_2_port, CK => clock, RB 
                           => resetn, Q => arx_state_reg_2_port);
   arx_o1_reg_reg_7 : DFERPQ1 port map( D => a_out_7_port, CEB => n175, CK => 
                           clock, RB => resetn, Q => data_out(7));
   arx_o1_reg_reg_0 : DFERPQ1 port map( D => a_out_0_port, CEB => n175, CK => 
                           clock, RB => resetn, Q => data_out(0));
   arx_o1_reg_reg_1 : DFERPQ1 port map( D => a_out_1_port, CEB => n175, CK => 
                           clock, RB => resetn, Q => data_out(1));
   arx_o1_reg_reg_2 : DFERPQ1 port map( D => a_out_2_port, CEB => n175, CK => 
                           clock, RB => resetn, Q => data_out(2));
   arx_o1_reg_reg_3 : DFERPQ1 port map( D => a_out_3_port, CEB => n175, CK => 
                           clock, RB => resetn, Q => data_out(3));
   arx_o1_reg_reg_4 : DFERPQ1 port map( D => a_out_4_port, CEB => n175, CK => 
                           clock, RB => resetn, Q => data_out(4));
   arx_o1_reg_reg_5 : DFERPQ1 port map( D => a_out_5_port, CEB => n175, CK => 
                           clock, RB => resetn, Q => data_out(5));
   arx_o1_reg_reg_6 : DFERPQ1 port map( D => a_out_6_port, CEB => n175, CK => 
                           clock, RB => resetn, Q => data_out(6));
   U205 : INVD1 port map( A => n99, Z => n178);
   U206 : NOR2D1 port map( A1 => m_in_l_0, A2 => m_in_l_4, Z => n99);
   U207 : NAN2D1 port map( A1 => n98, A2 => n99, Z => m2_in_l_3_port);
   U208 : NAN2M1D1 port map( A1 => m_in_l_4, A2 => n98, Z => m2_in_l_5_port);
   U209 : NAN2M1D1 port map( A1 => n67, A2 => n78, Z => state_0_port);
   U210 : INVD1 port map( A => n68, Z => n176);
   U211 : NAN2D1 port map( A1 => n63, A2 => n96, Z => m_in_l_4);
   U212 : AND2D1 port map( A1 => n100, A2 => n179, Z => n98);
   U213 : INVD1 port map( A => n77, Z => n179);
   U214 : NAN2D1 port map( A1 => n62, A2 => n78, Z => m_in_l_0);
   U215 : AND2D1 port map( A1 => n102, A2 => n96, Z => n101);
   U216 : NOR2M1D1 port map( A1 => n79, A2 => n67, Z => n102);
   U217 : NAN2D1 port map( A1 => n63, A2 => n100, Z => n67);
   U218 : NOR2D1 port map( A1 => n101, A2 => n199, Z => a_in_r_5_port);
   U219 : NOR2D1 port map( A1 => n102, A2 => n191, Z => a_in_l_6_port);
   U220 : NOR2D1 port map( A1 => n101, A2 => n198, Z => a_in_r_6_port);
   U221 : NOR2D1 port map( A1 => n102, A2 => n195, Z => a_in_l_2_port);
   U222 : NOR2D1 port map( A1 => n101, A2 => n202, Z => a_in_r_2_port);
   U223 : NOR2D1 port map( A1 => n102, A2 => n194, Z => a_in_l_3_port);
   U224 : NOR2D1 port map( A1 => n101, A2 => n201, Z => a_in_r_3_port);
   U225 : NOR2D1 port map( A1 => n102, A2 => n193, Z => a_in_l_4_port);
   U226 : NOR2D1 port map( A1 => n101, A2 => n200, Z => a_in_r_4_port);
   U227 : NOR2D1 port map( A1 => n102, A2 => n197, Z => a_in_l_0_port);
   U228 : NOR2D1 port map( A1 => n102, A2 => n196, Z => a_in_l_1_port);
   U229 : NOR2D1 port map( A1 => n101, A2 => n203, Z => a_in_r_1_port);
   U230 : NAN3D1 port map( A1 => n181, A2 => n182, A3 => n180, Z => n78);
   U231 : NOR2D1 port map( A1 => n101, A2 => n204, Z => a_in_r_0_port);
   U232 : NOR2D1 port map( A1 => n102, A2 => n192, Z => a_in_l_5_port);
   U233 : NOR2D1 port map( A1 => n101, A2 => n212, Z => a_in_r_14_port);
   U234 : NOR2M1D1 port map( A1 => n79, A2 => state_0_port, Z => n80);
   U235 : NAN3D1 port map( A1 => n62, A2 => n179, A3 => n80, Z => n64);
   U236 : NAN2D1 port map( A1 => n62, A2 => n96, Z => n68);
   U237 : OR3D1 port map( A1 => n77, A2 => state_0_port, A3 => n68, Z => n175);
   U238 : NAN4M1D1 port map( A1 => state_2_port, A2 => n79, A3 => n63, A4 => 
                           n62, Z => n97);
   U239 : NAN2D1 port map( A1 => n98, A2 => n96, Z => state_2_port);
   U240 : AND3D1 port map( A1 => n179, A2 => n78, A3 => n79, Z => n65);
   U241 : NAN3D1 port map( A1 => n62, A2 => n179, A3 => n63, Z => state_1_port)
                           ;
   U242 : NAN3D1 port map( A1 => arx_state_reg_0_port, A2 => n182, A3 => 
                           arx_state_reg_1_port, Z => n96);
   U243 : INVD1 port map( A => arx_state_reg_2_port, Z => n182);
   U244 : NOR3D1 port map( A1 => n180, A2 => arx_state_reg_1_port, A3 => n182, 
                           Z => n77);
   U245 : NAN3D1 port map( A1 => n181, A2 => n182, A3 => arx_state_reg_0_port, 
                           Z => n62);
   U246 : INVD1 port map( A => arx_state_reg_1_port, Z => n181);
   U247 : NAN3D1 port map( A1 => n180, A2 => n182, A3 => arx_state_reg_1_port, 
                           Z => n63);
   U248 : NOR2D1 port map( A1 => n101, A2 => n205, Z => a_in_r_7_port);
   U249 : NOR2D1 port map( A1 => n101, A2 => n206, Z => a_in_r_8_port);
   U250 : NOR2D1 port map( A1 => n101, A2 => n207, Z => a_in_r_9_port);
   U251 : NOR2D1 port map( A1 => n101, A2 => n208, Z => a_in_r_10_port);
   U252 : NOR2D1 port map( A1 => n101, A2 => n209, Z => a_in_r_11_port);
   U253 : NOR2D1 port map( A1 => n101, A2 => n210, Z => a_in_r_12_port);
   U254 : NOR2D1 port map( A1 => n101, A2 => n211, Z => a_in_r_13_port);
   U255 : INVD1 port map( A => arx_state_reg_0_port, Z => n180);
   U256 : NAN3D1 port map( A1 => n180, A2 => n181, A3 => arx_state_reg_2_port, 
                           Z => n100);
   U257 : NAN3D1 port map( A1 => arx_state_reg_1_port, A2 => n180, A3 => 
                           arx_state_reg_2_port, Z => n79);
   U258 : AND2D1 port map( A1 => N47, A2 => n178, Z => m_in_r_3_port);
   U259 : AND2D1 port map( A1 => N46, A2 => n178, Z => m_in_r_2_port);
   U260 : AND2D1 port map( A1 => N44, A2 => n178, Z => m_in_r_0_port);
   U261 : AND2D1 port map( A1 => N45, A2 => n178, Z => m_in_r_1_port);
   U262 : AND2D1 port map( A1 => N48, A2 => n178, Z => m_in_r_4_port);
   U263 : AND2D1 port map( A1 => N50, A2 => n178, Z => m_in_r_6_port);
   U264 : AND2D1 port map( A1 => N49, A2 => n178, Z => m_in_r_5_port);
   U265 : AND2D1 port map( A1 => N51, A2 => n178, Z => m_in_r_7_port);
   U266 : INVD1 port map( A => arx_r2_reg_1_port, Z => n203);
   U267 : INVD1 port map( A => arx_r1_reg_1_port, Z => n196);
   U268 : INVD1 port map( A => arx_r1_reg_0_port, Z => n197);
   U269 : INVD1 port map( A => arx_r2_reg_0_port, Z => n204);
   U270 : INVD1 port map( A => arx_r1_reg_2_port, Z => n195);
   U271 : INVD1 port map( A => arx_r2_reg_2_port, Z => n202);
   U272 : INVD1 port map( A => arx_r1_reg_3_port, Z => n194);
   U273 : INVD1 port map( A => arx_r2_reg_3_port, Z => n201);
   U274 : INVD1 port map( A => arx_r1_reg_4_port, Z => n193);
   U275 : INVD1 port map( A => arx_r2_reg_4_port, Z => n200);
   U276 : INVD1 port map( A => arx_r1_reg_5_port, Z => n192);
   U277 : INVD1 port map( A => arx_r2_reg_5_port, Z => n199);
   U278 : INVD1 port map( A => arx_r2_reg_6_port, Z => n198);
   U279 : INVD1 port map( A => arx_r1_reg_6_port, Z => n191);
   U280 : INVD1 port map( A => arx_r1_reg_7_port, Z => n190);
   U281 : INVD1 port map( A => arx_r2_reg_7_port, Z => n205);
   U282 : INVD1 port map( A => arx_r1_reg_8_port, Z => n189);
   U283 : INVD1 port map( A => arx_r2_reg_8_port, Z => n206);
   U284 : INVD1 port map( A => arx_r1_reg_9_port, Z => n188);
   U285 : INVD1 port map( A => arx_r2_reg_9_port, Z => n207);
   U286 : INVD1 port map( A => arx_r1_reg_10_port, Z => n187);
   U287 : INVD1 port map( A => arx_r2_reg_10_port, Z => n208);
   U288 : INVD1 port map( A => arx_r1_reg_11_port, Z => n186);
   U289 : INVD1 port map( A => arx_r2_reg_11_port, Z => n209);
   U290 : INVD1 port map( A => arx_r1_reg_12_port, Z => n185);
   U291 : INVD1 port map( A => arx_r2_reg_12_port, Z => n210);
   U292 : INVD1 port map( A => arx_r1_reg_13_port, Z => n184);
   U293 : INVD1 port map( A => arx_r2_reg_13_port, Z => n211);
   U294 : INVD1 port map( A => arx_r1_reg_14_port, Z => n183);
   U295 : INVD1 port map( A => arx_r2_reg_14_port, Z => n212);
   U296 : TIELO port map( Z => net1366);
   U297 : EXOR2D1 port map( A1 => N152, A2 => add_416_C204_rn_carry_7_port, Z 
                           => a_out_7_port);
   U298 : AND2D1 port map( A1 => add_416_C204_rn_carry_6_port, A2 => N151, Z =>
                           add_416_C204_rn_carry_7_port);
   U299 : EXOR2D1 port map( A1 => N151, A2 => add_416_C204_rn_carry_6_port, Z 
                           => a_out_6_port);
   U300 : AND2D1 port map( A1 => add_416_C204_rn_carry_5_port, A2 => N150, Z =>
                           add_416_C204_rn_carry_6_port);
   U301 : EXOR2D1 port map( A1 => N150, A2 => add_416_C204_rn_carry_5_port, Z 
                           => a_out_5_port);
   U302 : AND2D1 port map( A1 => add_416_C204_rn_carry_4_port, A2 => N149, Z =>
                           add_416_C204_rn_carry_5_port);
   U303 : EXOR2D1 port map( A1 => N149, A2 => add_416_C204_rn_carry_4_port, Z 
                           => a_out_4_port);
   U304 : AND2D1 port map( A1 => add_416_C204_rn_carry_3_port, A2 => N148, Z =>
                           add_416_C204_rn_carry_4_port);
   U305 : EXOR2D1 port map( A1 => N148, A2 => add_416_C204_rn_carry_3_port, Z 
                           => a_out_3_port);
   U306 : AND2D1 port map( A1 => add_416_C204_rn_carry_2_port, A2 => N147, Z =>
                           add_416_C204_rn_carry_3_port);
   U307 : EXOR2D1 port map( A1 => N147, A2 => add_416_C204_rn_carry_2_port, Z 
                           => a_out_2_port);
   U308 : AND2D1 port map( A1 => add_416_C204_rn_carry_1_port, A2 => N146, Z =>
                           add_416_C204_rn_carry_2_port);
   U309 : EXOR2D1 port map( A1 => N146, A2 => add_416_C204_rn_carry_1_port, Z 
                           => a_out_1_port);
   U310 : AND2D1 port map( A1 => N145, A2 => N144, Z => 
                           add_416_C204_rn_carry_1_port);
   U311 : EXOR2D1 port map( A1 => N144, A2 => N145, Z => a_out_0_port);
   U312 : NOR2D1 port map( A1 => arx_state_reg_1_port, A2 => n182, Z => n177);
   U313 : AO22D1 port map( A1 => N52, A2 => n182, B1 => N44, B2 => n177, Z => 
                           m2_in_r_0_port);
   U314 : AO22D1 port map( A1 => N53, A2 => n182, B1 => N45, B2 => n177, Z => 
                           m2_in_r_1_port);
   U315 : AO22D1 port map( A1 => N54, A2 => n182, B1 => N46, B2 => n177, Z => 
                           m2_in_r_2_port);
   U316 : AO22D1 port map( A1 => N55, A2 => n182, B1 => N47, B2 => n177, Z => 
                           m2_in_r_3_port);
   U317 : AO22D1 port map( A1 => N56, A2 => n182, B1 => N48, B2 => n177, Z => 
                           m2_in_r_4_port);
   U318 : AO22D1 port map( A1 => N57, A2 => n182, B1 => N49, B2 => n177, Z => 
                           m2_in_r_5_port);
   U319 : AO22D1 port map( A1 => N58, A2 => n182, B1 => N50, B2 => n177, Z => 
                           m2_in_r_6_port);
   U320 : AO22D1 port map( A1 => N59, A2 => n182, B1 => N51, B2 => n177, Z => 
                           m2_in_r_7_port);
   add_204_U10 : OAI211D1 port map( A1 => a_in_l_1_port, A2 => a_in_r_1_port, B
                           => a_in_l_0_port, C => a_in_r_0_port, Z => 
                           add_204_n9);
   add_204_U9 : OAI21M20D1 port map( A1 => a_in_l_1_port, A2 => a_in_r_1_port, 
                           B => add_204_n9, Z => add_204_n7);
   add_204_U8 : OAI21D1 port map( A1 => a_in_l_2_port, A2 => add_204_n7, B => 
                           a_in_r_2_port, Z => add_204_n8);
   add_204_U7 : OAI21M20D1 port map( A1 => add_204_n7, A2 => a_in_l_2_port, B 
                           => add_204_n8, Z => add_204_n5);
   add_204_U6 : OAI21D1 port map( A1 => a_in_l_3_port, A2 => add_204_n5, B => 
                           a_in_r_3_port, Z => add_204_n6);
   add_204_U5 : OAI21M20D1 port map( A1 => add_204_n5, A2 => a_in_l_3_port, B 
                           => add_204_n6, Z => add_204_n3);
   add_204_U4 : OAI21D1 port map( A1 => a_in_l_4_port, A2 => add_204_n3, B => 
                           a_in_r_4_port, Z => add_204_n4);
   add_204_U3 : OAI21M20D1 port map( A1 => add_204_n3, A2 => a_in_l_4_port, B 
                           => add_204_n4, Z => add_204_n1);
   add_204_U2 : OAI21D1 port map( A1 => a_in_l_5_port, A2 => add_204_n1, B => 
                           a_in_r_5_port, Z => add_204_n2);
   add_204_U1 : OAI21M20D1 port map( A1 => add_204_n1, A2 => a_in_l_5_port, B 
                           => add_204_n2, Z => add_204_carry_6_port);
   add_204_U1_14 : EXOR3D1 port map( A1 => a_in_l_14_port, A2 => a_in_r_14_port
                           , A3 => add_204_carry_14_port, Z => N152);
   add_204_U1_6 : ADFULD1 port map( A => a_in_l_6_port, B => a_in_r_6_port, CI 
                           => add_204_carry_6_port, CO => add_204_carry_7_port,
                           S => N144);
   add_204_U1_7 : ADFULD1 port map( A => a_in_l_7_port, B => a_in_r_7_port, CI 
                           => add_204_carry_7_port, CO => add_204_carry_8_port,
                           S => N145);
   add_204_U1_8 : ADFULD1 port map( A => a_in_l_8_port, B => a_in_r_8_port, CI 
                           => add_204_carry_8_port, CO => add_204_carry_9_port,
                           S => N146);
   add_204_U1_9 : ADFULD1 port map( A => a_in_l_9_port, B => a_in_r_9_port, CI 
                           => add_204_carry_9_port, CO => add_204_carry_10_port
                           , S => N147);
   add_204_U1_10 : ADFULD1 port map( A => a_in_l_10_port, B => a_in_r_10_port, 
                           CI => add_204_carry_10_port, CO => 
                           add_204_carry_11_port, S => N148);
   add_204_U1_11 : ADFULD1 port map( A => a_in_l_11_port, B => a_in_r_11_port, 
                           CI => add_204_carry_11_port, CO => 
                           add_204_carry_12_port, S => N149);
   add_204_U1_12 : ADFULD1 port map( A => a_in_l_12_port, B => a_in_r_12_port, 
                           CI => add_204_carry_12_port, CO => 
                           add_204_carry_13_port, S => N150);
   add_204_U1_13 : ADFULD1 port map( A => a_in_l_13_port, B => a_in_r_13_port, 
                           CI => add_204_carry_13_port, CO => 
                           add_204_carry_14_port, S => N151);
   mult_203_U232 : EXOR2D1 port map( A1 => m_in_l_0, A2 => m2_in_l_5_port, Z =>
                           mult_203_n208);
   mult_203_U231 : EXOR2D1 port map( A1 => m2_in_r_7_port, A2 => m_in_l_0, Z =>
                           mult_203_n209);
   mult_203_U230 : EXNOR2D1 port map( A1 => m2_in_r_6_port, A2 => mult_203_n203
                           , Z => mult_203_n237);
   mult_203_U229 : EXNOR2D1 port map( A1 => m2_in_r_7_port, A2 => 
                           m2_in_l_5_port, Z => mult_203_n231);
   mult_203_U228 : EXOR2D1 port map( A1 => m2_in_r_6_port, A2 => mult_203_n206,
                           Z => mult_203_n230);
   mult_203_U227 : EXOR2D1 port map( A1 => m2_in_r_6_port, A2 => mult_203_n205,
                           Z => mult_203_n240);
   mult_203_U226 : EXOR2D1 port map( A1 => m2_in_l_3_port, A2 => m_in_l_0, Z =>
                           mult_203_n241);
   mult_203_U225 : EXOR2D1 port map( A1 => m2_in_r_2_port, A2 => mult_203_n203,
                           Z => mult_203_n234);
   mult_203_U224 : EXOR2D1 port map( A1 => m2_in_r_1_port, A2 => mult_203_n203,
                           Z => mult_203_n232);
   mult_203_U223 : EXOR2D1 port map( A1 => m2_in_r_5_port, A2 => mult_203_n205,
                           Z => mult_203_n223);
   mult_203_U222 : OR2D1 port map( A1 => mult_203_n238, A2 => mult_203_n239, Z 
                           => mult_203_n37);
   mult_203_U221 : EXNOR2D1 port map( A1 => mult_203_n238, A2 => mult_203_n239,
                           Z => mult_203_n38);
   mult_203_U220 : OAI21D1 port map( A1 => m2_in_r_0_port, A2 => mult_203_n203,
                           B => mult_203_n211, Z => mult_203_n60);
   mult_203_U219 : EXOR2D1 port map( A1 => m2_in_r_5_port, A2 => mult_203_n203,
                           Z => mult_203_n236);
   mult_203_U218 : EXOR2D1 port map( A1 => m2_in_r_4_port, A2 => mult_203_n203,
                           Z => mult_203_n235);
   mult_203_U217 : EXOR2D1 port map( A1 => m2_in_r_3_port, A2 => mult_203_n203,
                           Z => mult_203_n233);
   mult_203_U216 : NOR2D1 port map( A1 => mult_203_n201, A2 => mult_203_n200, Z
                           => mult_203_n68);
   mult_203_U215 : EXOR2D1 port map( A1 => m2_in_r_5_port, A2 => mult_203_n206,
                           Z => mult_203_n229);
   mult_203_U214 : EXOR2D1 port map( A1 => m2_in_r_4_port, A2 => mult_203_n206,
                           Z => mult_203_n228);
   mult_203_U213 : EXOR2D1 port map( A1 => m2_in_r_3_port, A2 => mult_203_n206,
                           Z => mult_203_n227);
   mult_203_U212 : EXOR2D1 port map( A1 => m2_in_r_2_port, A2 => mult_203_n206,
                           Z => mult_203_n226);
   mult_203_U211 : EXOR2D1 port map( A1 => m2_in_r_1_port, A2 => mult_203_n206,
                           Z => mult_203_n225);
   mult_203_U210 : NOR2D1 port map( A1 => mult_203_n224, A2 => mult_203_n200, Z
                           => mult_203_n76);
   mult_203_U209 : EXOR2D1 port map( A1 => m2_in_r_4_port, A2 => mult_203_n205,
                           Z => mult_203_n222);
   mult_203_U208 : EXOR2D1 port map( A1 => m2_in_r_3_port, A2 => mult_203_n205,
                           Z => mult_203_n221);
   mult_203_U207 : EXOR2D1 port map( A1 => m2_in_r_2_port, A2 => mult_203_n205,
                           Z => mult_203_n220);
   mult_203_U206 : EXOR2D1 port map( A1 => m2_in_r_1_port, A2 => mult_203_n205,
                           Z => mult_203_n218);
   mult_203_U205 : EXOR2D1 port map( A1 => mult_203_n205, A2 => m2_in_r_0_port,
                           Z => mult_203_n219);
   mult_203_U204 : EXNOR2D1 port map( A1 => m2_in_r_7_port, A2 => m_in_l_0, Z 
                           => mult_203_n217);
   mult_203_U203 : AO21D1 port map( A1 => mult_203_n205, A2 => mult_203_n211, B
                           => mult_203_n217, Z => mult_203_n85);
   mult_203_U202 : EXOR2D1 port map( A1 => m2_in_r_6_port, A2 => mult_203_n203,
                           Z => mult_203_n216);
   mult_203_U201 : OAI22D1 port map( A1 => mult_203_n217, A2 => mult_203_n205, 
                           B1 => mult_203_n216, B2 => mult_203_n211, Z => 
                           mult_203_n86);
   mult_203_U200 : EXOR2D1 port map( A1 => m2_in_r_5_port, A2 => mult_203_n203,
                           Z => mult_203_n215);
   mult_203_U199 : OAI22D1 port map( A1 => mult_203_n216, A2 => mult_203_n205, 
                           B1 => mult_203_n215, B2 => mult_203_n211, Z => 
                           mult_203_n87);
   mult_203_U198 : EXOR2D1 port map( A1 => m2_in_r_4_port, A2 => mult_203_n203,
                           Z => mult_203_n214);
   mult_203_U197 : OAI22D1 port map( A1 => mult_203_n215, A2 => mult_203_n205, 
                           B1 => mult_203_n214, B2 => mult_203_n211, Z => 
                           mult_203_n88);
   mult_203_U196 : EXOR2D1 port map( A1 => m2_in_r_3_port, A2 => mult_203_n203,
                           Z => mult_203_n213);
   mult_203_U195 : OAI22D1 port map( A1 => mult_203_n214, A2 => mult_203_n205, 
                           B1 => mult_203_n213, B2 => mult_203_n211, Z => 
                           mult_203_n89);
   mult_203_U194 : EXOR2D1 port map( A1 => m2_in_r_2_port, A2 => mult_203_n203,
                           Z => mult_203_n212);
   mult_203_U193 : OAI22D1 port map( A1 => mult_203_n213, A2 => mult_203_n205, 
                           B1 => mult_203_n212, B2 => mult_203_n211, Z => 
                           mult_203_n90);
   mult_203_U192 : EXOR2D1 port map( A1 => m2_in_r_1_port, A2 => mult_203_n203,
                           Z => mult_203_n210);
   mult_203_U191 : OAI22D1 port map( A1 => mult_203_n212, A2 => mult_203_n205, 
                           B1 => mult_203_n210, B2 => mult_203_n211, Z => 
                           mult_203_n91);
   mult_203_U190 : OAI22D1 port map( A1 => mult_203_n210, A2 => mult_203_n205, 
                           B1 => m2_in_r_0_port, B2 => mult_203_n211, Z => 
                           mult_203_n92);
   mult_203_U189 : NOR2D1 port map( A1 => mult_203_n205, A2 => mult_203_n200, Z
                           => m2_out_0_port);
   mult_203_U188 : EXNOR3D1 port map( A1 => mult_203_n2, A2 => mult_203_n16, A3
                           => mult_203_n207, Z => m2_out_14_port);
   mult_203_U187 : EXOR2D1 port map( A1 => mult_203_n91, A2 => mult_203_n14, Z 
                           => m2_out_2_port);
   mult_203_U186 : INVD1 port map( A => mult_203_n21, Z => mult_203_n197);
   mult_203_U185 : NOR2D1 port map( A1 => mult_203_n201, A2 => mult_203_n236, Z
                           => mult_203_n63);
   mult_203_U184 : NOR2D1 port map( A1 => mult_203_n224, A2 => mult_203_n230, Z
                           => mult_203_n70);
   mult_203_U183 : NOR2D1 port map( A1 => mult_203_n201, A2 => mult_203_n235, Z
                           => mult_203_n64);
   mult_203_U182 : EXOR2D1 port map( A1 => m2_in_r_7_port, A2 => m2_in_l_3_port
                           , Z => mult_203_n195);
   mult_203_U181 : NOR2D1 port map( A1 => mult_203_n240, A2 => mult_203_n202, Z
                           => mult_203_n31);
   mult_203_U180 : NOR2D1 port map( A1 => mult_203_n201, A2 => mult_203_n234, Z
                           => mult_203_n238);
   mult_203_U179 : NOR2D1 port map( A1 => mult_203_n223, A2 => mult_203_n202, Z
                           => mult_203_n239);
   mult_203_U178 : INVD1 port map( A => m2_in_r_0_port, Z => mult_203_n200);
   mult_203_U177 : NOR2D1 port map( A1 => mult_203_n224, A2 => mult_203_n228, Z
                           => mult_203_n72);
   mult_203_U176 : NOR3D1 port map( A1 => mult_203_n201, A2 => mult_203_n203, 
                           A3 => m2_in_r_0_port, Z => mult_203_n57);
   mult_203_U175 : NOR2D1 port map( A1 => mult_203_n224, A2 => mult_203_n226, Z
                           => mult_203_n74);
   mult_203_U174 : NOR3D1 port map( A1 => mult_203_n224, A2 => mult_203_n206, 
                           A3 => m2_in_r_0_port, Z => mult_203_n58);
   mult_203_U173 : NOR2D1 port map( A1 => mult_203_n224, A2 => mult_203_n225, Z
                           => mult_203_n75);
   mult_203_U172 : NOR2D1 port map( A1 => mult_203_n220, A2 => mult_203_n202, Z
                           => mult_203_n81);
   mult_203_U171 : NOR2D1 port map( A1 => mult_203_n219, A2 => mult_203_n202, Z
                           => mult_203_n83);
   mult_203_U170 : NAN2D1 port map( A1 => mult_203_n208, A2 => mult_203_n209, Z
                           => mult_203_n16);
   mult_203_U169 : INVD1 port map( A => mult_203_n231, Z => mult_203_n196);
   mult_203_U168 : INVD1 port map( A => mult_203_n237, Z => mult_203_n199);
   mult_203_U167 : NAN2D1 port map( A1 => mult_203_n204, A2 => mult_203_n196, Z
                           => mult_203_n69);
   mult_203_U166 : NOR2D1 port map( A1 => mult_203_n201, A2 => mult_203_n199, Z
                           => mult_203_n62);
   mult_203_U165 : NOR2D1 port map( A1 => mult_203_n224, A2 => mult_203_n231, Z
                           => mult_203_n21);
   mult_203_U164 : INVD1 port map( A => mult_203_n31, Z => mult_203_n198);
   mult_203_U163 : NOR2D1 port map( A1 => mult_203_n224, A2 => mult_203_n229, Z
                           => mult_203_n71);
   mult_203_U162 : NOR2D1 port map( A1 => mult_203_n201, A2 => mult_203_n233, Z
                           => mult_203_n65);
   mult_203_U161 : NOR2D1 port map( A1 => mult_203_n222, A2 => mult_203_n202, Z
                           => mult_203_n79);
   mult_203_U160 : NOR2D1 port map( A1 => mult_203_n201, A2 => mult_203_n232, Z
                           => mult_203_n67);
   mult_203_U159 : NOR2D1 port map( A1 => mult_203_n224, A2 => mult_203_n227, Z
                           => mult_203_n73);
   mult_203_U158 : INVD1 port map( A => m_in_l_0, Z => mult_203_n203);
   mult_203_U157 : NOR2D1 port map( A1 => mult_203_n221, A2 => mult_203_n202, Z
                           => mult_203_n80);
   mult_203_U156 : NAN2D1 port map( A1 => m_in_l_0, A2 => mult_203_n205, Z => 
                           mult_203_n211);
   mult_203_U155 : NOR2D1 port map( A1 => mult_203_n218, A2 => mult_203_n202, Z
                           => mult_203_n82);
   mult_203_U154 : NOR2D1 port map( A1 => mult_203_n205, A2 => mult_203_n202, Z
                           => mult_203_n59);
   mult_203_U153 : NAN2D1 port map( A1 => mult_203_n208, A2 => mult_203_n209, Z
                           => mult_203_n207);
   mult_203_U152 : INVD1 port map( A => m2_in_l_5_port, Z => mult_203_n206);
   mult_203_U151 : INVD1 port map( A => mult_203_n208, Z => mult_203_n201);
   mult_203_U150 : INVD1 port map( A => m2_in_l_3_port, Z => mult_203_n205);
   mult_203_U149 : EXOR2D1 port map( A1 => m2_in_l_5_port, A2 => mult_203_n205,
                           Z => mult_203_n224);
   mult_203_U148 : INVD1 port map( A => mult_203_n241, Z => mult_203_n202);
   mult_203_U147 : INVD1 port map( A => mult_203_n224, Z => mult_203_n204);
   mult_203_U146 : NAN2D1 port map( A1 => mult_203_n241, A2 => mult_203_n195, Z
                           => mult_203_n77);
   mult_203_U145 : AND2D1 port map( A1 => mult_203_n14, A2 => mult_203_n91, Z 
                           => mult_203_n194);
   mult_203_U37 : ADHALFDL port map( A => mult_203_n83, B => mult_203_n90, CO 
                           => mult_203_n55, S => mult_203_n56);
   mult_203_U36 : ADFULD1 port map( A => mult_203_n89, B => mult_203_n76, CI =>
                           mult_203_n82, CO => mult_203_n53, S => mult_203_n54)
                           ;
   mult_203_U35 : ADHALFDL port map( A => mult_203_n58, B => mult_203_n88, CO 
                           => mult_203_n51, S => mult_203_n52);
   mult_203_U34 : ADFULD1 port map( A => mult_203_n75, B => mult_203_n81, CI =>
                           mult_203_n52, CO => mult_203_n49, S => mult_203_n50)
                           ;
   mult_203_U33 : ADFULD1 port map( A => mult_203_n87, B => mult_203_n68, CI =>
                           mult_203_n80, CO => mult_203_n47, S => mult_203_n48)
                           ;
   mult_203_U32 : ADFULD1 port map( A => mult_203_n51, B => mult_203_n74, CI =>
                           mult_203_n48, CO => mult_203_n45, S => mult_203_n46)
                           ;
   mult_203_U31 : ADHALFDL port map( A => mult_203_n57, B => mult_203_n86, CO 
                           => mult_203_n43, S => mult_203_n44);
   mult_203_U30 : ADFULD1 port map( A => mult_203_n67, B => mult_203_n79, CI =>
                           mult_203_n73, CO => mult_203_n41, S => mult_203_n42)
                           ;
   mult_203_U29 : ADFULD1 port map( A => mult_203_n47, B => mult_203_n44, CI =>
                           mult_203_n42, CO => mult_203_n39, S => mult_203_n40)
                           ;
   mult_203_U26 : ADFULD1 port map( A => mult_203_n85, B => mult_203_n72, CI =>
                           mult_203_n43, CO => mult_203_n35, S => mult_203_n36)
                           ;
   mult_203_U25 : ADFULD1 port map( A => mult_203_n41, B => mult_203_n38, CI =>
                           mult_203_n36, CO => mult_203_n33, S => mult_203_n34)
                           ;
   mult_203_U23 : ADFULD1 port map( A => mult_203_n65, B => mult_203_n71, CI =>
                           mult_203_n198, CO => mult_203_n29, S => mult_203_n30
                           );
   mult_203_U22 : ADFULD1 port map( A => mult_203_n35, B => mult_203_n37, CI =>
                           mult_203_n30, CO => mult_203_n27, S => mult_203_n28)
                           ;
   mult_203_U21 : ADFULD1 port map( A => mult_203_n70, B => mult_203_n31, CI =>
                           mult_203_n64, CO => mult_203_n25, S => mult_203_n26)
                           ;
   mult_203_U20 : ADFULD1 port map( A => mult_203_n29, B => mult_203_n77, CI =>
                           mult_203_n26, CO => mult_203_n23, S => mult_203_n24)
                           ;
   mult_203_U18 : ADFULD1 port map( A => mult_203_n197, B => mult_203_n63, CI 
                           => mult_203_n25, CO => mult_203_n19, S => 
                           mult_203_n20);
   mult_203_U17 : ADFULD1 port map( A => mult_203_n62, B => mult_203_n21, CI =>
                           mult_203_n69, CO => mult_203_n17, S => mult_203_n18)
                           ;
   mult_203_U15 : ADHALFDL port map( A => mult_203_n92, B => mult_203_n60, CO 
                           => mult_203_n14, S => m2_out_1_port);
   mult_203_U13 : ADFULD1 port map( A => mult_203_n56, B => mult_203_n59, CI =>
                           mult_203_n194, CO => mult_203_n12, S => 
                           m2_out_3_port);
   mult_203_U12 : ADFULD1 port map( A => mult_203_n54, B => mult_203_n55, CI =>
                           mult_203_n12, CO => mult_203_n11, S => m2_out_4_port
                           );
   mult_203_U11 : ADFULD1 port map( A => mult_203_n50, B => mult_203_n53, CI =>
                           mult_203_n11, CO => mult_203_n10, S => m2_out_5_port
                           );
   mult_203_U10 : ADFULD1 port map( A => mult_203_n46, B => mult_203_n49, CI =>
                           mult_203_n10, CO => mult_203_n9, S => m2_out_6_port)
                           ;
   mult_203_U9 : ADFULD1 port map( A => mult_203_n40, B => mult_203_n45, CI => 
                           mult_203_n9, CO => mult_203_n8, S => m2_out_7_port);
   mult_203_U8 : ADFULD1 port map( A => mult_203_n34, B => mult_203_n39, CI => 
                           mult_203_n8, CO => mult_203_n7, S => m2_out_8_port);
   mult_203_U7 : ADFULD1 port map( A => mult_203_n28, B => mult_203_n33, CI => 
                           mult_203_n7, CO => mult_203_n6, S => m2_out_9_port);
   mult_203_U6 : ADFULD1 port map( A => mult_203_n24, B => mult_203_n27, CI => 
                           mult_203_n6, CO => mult_203_n5, S => m2_out_10_port)
                           ;
   mult_203_U5 : ADFULD1 port map( A => mult_203_n20, B => mult_203_n23, CI => 
                           mult_203_n5, CO => mult_203_n4, S => m2_out_11_port)
                           ;
   mult_203_U4 : ADFULD1 port map( A => mult_203_n19, B => mult_203_n18, CI => 
                           mult_203_n4, CO => mult_203_n3, S => m2_out_12_port)
                           ;
   mult_203_U3 : ADFULD1 port map( A => mult_203_n17, B => mult_203_n16, CI => 
                           mult_203_n3, CO => mult_203_n2, S => m2_out_13_port)
                           ;
   mult_202_U172 : NOR2D1 port map( A1 => mult_202_n177, A2 => mult_202_n178, Z
                           => mult_202_n100);
   mult_202_U171 : NAN2D1 port map( A1 => n178, A2 => m_in_r_7_port, Z => 
                           mult_202_n101);
   mult_202_U170 : NOR2D1 port map( A1 => mult_202_n169, A2 => mult_202_n176, Z
                           => mult_202_n102);
   mult_202_U169 : NOR2D1 port map( A1 => mult_202_n170, A2 => mult_202_n176, Z
                           => mult_202_n103);
   mult_202_U168 : NOR2D1 port map( A1 => mult_202_n171, A2 => mult_202_n176, Z
                           => mult_202_n104);
   mult_202_U167 : NOR2D1 port map( A1 => mult_202_n172, A2 => mult_202_n176, Z
                           => mult_202_n105);
   mult_202_U166 : NOR2D1 port map( A1 => mult_202_n173, A2 => mult_202_n176, Z
                           => mult_202_n106);
   mult_202_U165 : NOR2D1 port map( A1 => mult_202_n174, A2 => mult_202_n176, Z
                           => mult_202_n107);
   mult_202_U164 : NOR2D1 port map( A1 => mult_202_n177, A2 => mult_202_n176, Z
                           => mult_202_n108);
   mult_202_U163 : NAN2D1 port map( A1 => m_in_l_0, A2 => m_in_r_7_port, Z => 
                           mult_202_n109);
   mult_202_U162 : NOR2D1 port map( A1 => mult_202_n175, A2 => mult_202_n169, Z
                           => mult_202_n110);
   mult_202_U161 : NOR2D1 port map( A1 => mult_202_n175, A2 => mult_202_n170, Z
                           => mult_202_n111);
   mult_202_U160 : NOR2D1 port map( A1 => mult_202_n175, A2 => mult_202_n171, Z
                           => mult_202_n112);
   mult_202_U159 : NOR2D1 port map( A1 => mult_202_n175, A2 => mult_202_n172, Z
                           => mult_202_n113);
   mult_202_U158 : NOR2D1 port map( A1 => mult_202_n175, A2 => mult_202_n173, Z
                           => mult_202_n114);
   mult_202_U157 : NOR2D1 port map( A1 => mult_202_n175, A2 => mult_202_n174, Z
                           => mult_202_n115);
   mult_202_U156 : NAN2D1 port map( A1 => m_in_l_0, A2 => m_in_r_6_port, Z => 
                           mult_202_n20);
   mult_202_U155 : NAN2D1 port map( A1 => m_in_r_6_port, A2 => m_in_l_4, Z => 
                           mult_202_n38);
   mult_202_U154 : NAN2D1 port map( A1 => m_in_r_5_port, A2 => m_in_l_4, Z => 
                           mult_202_n181);
   mult_202_U153 : NAN2D1 port map( A1 => m_in_l_0, A2 => m_in_r_2_port, Z => 
                           mult_202_n180);
   mult_202_U152 : NAN2D1 port map( A1 => mult_202_n181, A2 => mult_202_n180, Z
                           => mult_202_n45);
   mult_202_U151 : EXNOR2D1 port map( A1 => mult_202_n180, A2 => mult_202_n181,
                           Z => mult_202_n46);
   mult_202_U150 : NAN2D1 port map( A1 => m_in_r_6_port, A2 => m_in_l_4, Z => 
                           mult_202_n72);
   mult_202_U149 : NAN2D1 port map( A1 => m_in_r_5_port, A2 => m_in_l_4, Z => 
                           mult_202_n73);
   mult_202_U148 : NAN2D1 port map( A1 => m_in_r_4_port, A2 => m_in_l_4, Z => 
                           mult_202_n74);
   mult_202_U147 : NAN2D1 port map( A1 => m_in_r_3_port, A2 => m_in_l_4, Z => 
                           mult_202_n75);
   mult_202_U146 : NAN2D1 port map( A1 => m_in_r_2_port, A2 => m_in_l_4, Z => 
                           mult_202_n76);
   mult_202_U145 : NAN2D1 port map( A1 => m_in_r_1_port, A2 => m_in_l_4, Z => 
                           mult_202_n77);
   mult_202_U144 : NAN2D1 port map( A1 => m_in_r_0_port, A2 => m_in_l_4, Z => 
                           mult_202_n78);
   mult_202_U143 : NAN2D1 port map( A1 => m_in_l_0, A2 => m_in_r_7_port, Z => 
                           mult_202_n79);
   mult_202_U142 : NOR2D1 port map( A1 => mult_202_n170, A2 => mult_202_n175, Z
                           => mult_202_n80);
   mult_202_U141 : NOR2D1 port map( A1 => mult_202_n171, A2 => mult_202_n175, Z
                           => mult_202_n81);
   mult_202_U140 : NOR2D1 port map( A1 => mult_202_n172, A2 => mult_202_n175, Z
                           => mult_202_n82);
   mult_202_U139 : NOR2D1 port map( A1 => mult_202_n174, A2 => mult_202_n175, Z
                           => mult_202_n84);
   mult_202_U138 : NOR2D1 port map( A1 => mult_202_n177, A2 => mult_202_n175, Z
                           => mult_202_n85);
   mult_202_U137 : NAN2D1 port map( A1 => m_in_l_4, A2 => m_in_r_7_port, Z => 
                           mult_202_n86);
   mult_202_U136 : NOR2D1 port map( A1 => mult_202_n178, A2 => mult_202_n169, Z
                           => mult_202_n87);
   mult_202_U135 : NOR2D1 port map( A1 => mult_202_n178, A2 => mult_202_n170, Z
                           => mult_202_n88);
   mult_202_U134 : NOR2D1 port map( A1 => mult_202_n171, A2 => mult_202_n178, Z
                           => mult_202_n89);
   mult_202_U133 : NOR2D1 port map( A1 => mult_202_n172, A2 => mult_202_n178, Z
                           => mult_202_n90);
   mult_202_U132 : NOR2D1 port map( A1 => mult_202_n173, A2 => mult_202_n178, Z
                           => mult_202_n91);
   mult_202_U131 : NOR2D1 port map( A1 => mult_202_n174, A2 => mult_202_n178, Z
                           => mult_202_n92);
   mult_202_U130 : NOR2D1 port map( A1 => mult_202_n177, A2 => mult_202_n178, Z
                           => mult_202_n93);
   mult_202_U129 : NAN2D1 port map( A1 => m_in_l_4, A2 => m_in_r_7_port, Z => 
                           mult_202_n94);
   mult_202_U128 : NOR2D1 port map( A1 => mult_202_n178, A2 => mult_202_n171, Z
                           => mult_202_n96);
   mult_202_U127 : NOR2D1 port map( A1 => mult_202_n178, A2 => mult_202_n172, Z
                           => mult_202_n97);
   mult_202_U126 : NOR2D1 port map( A1 => mult_202_n178, A2 => mult_202_n173, Z
                           => mult_202_n98);
   mult_202_U125 : NOR2D1 port map( A1 => mult_202_n178, A2 => mult_202_n174, Z
                           => mult_202_n99);
   mult_202_U124 : NOR2D1 port map( A1 => mult_202_n175, A2 => mult_202_n177, Z
                           => m_out_0_port);
   mult_202_U123 : AND2D1 port map( A1 => m_in_l_4, A2 => m_in_r_7_port, Z => 
                           mult_202_n179);
   mult_202_U122 : EXOR3D1 port map( A1 => mult_202_n2, A2 => mult_202_n15, A3 
                           => mult_202_n179, Z => m_out_14_port);
   mult_202_U121 : INVD1 port map( A => mult_202_n20, Z => mult_202_n168);
   mult_202_U120 : INVD1 port map( A => mult_202_n38, Z => mult_202_n167);
   mult_202_U119 : INVD1 port map( A => m_in_r_5_port, Z => mult_202_n170);
   mult_202_U118 : INVD1 port map( A => m_in_r_6_port, Z => mult_202_n169);
   mult_202_U117 : INVD1 port map( A => m_in_r_4_port, Z => mult_202_n171);
   mult_202_U116 : INVD1 port map( A => m_in_r_1_port, Z => mult_202_n174);
   mult_202_U115 : INVD1 port map( A => m_in_r_0_port, Z => mult_202_n177);
   mult_202_U114 : INVD1 port map( A => m_in_r_2_port, Z => mult_202_n173);
   mult_202_U113 : INVD1 port map( A => m_in_r_3_port, Z => mult_202_n172);
   mult_202_U112 : INVD1 port map( A => m_in_l_4, Z => mult_202_n178);
   mult_202_U111 : INVD1 port map( A => m_in_l_0, Z => mult_202_n175);
   mult_202_U110 : INVD1 port map( A => n178, Z => mult_202_n176);
   mult_202_U44 : ADHALFDL port map( A => mult_202_n106, B => mult_202_n113, CO
                           => mult_202_n69, S => mult_202_n70);
   mult_202_U43 : ADHALFDL port map( A => mult_202_n93, B => mult_202_n99, CO 
                           => mult_202_n67, S => mult_202_n68);
   mult_202_U42 : ADFULD1 port map( A => mult_202_n105, B => mult_202_n112, CI 
                           => mult_202_n69, CO => mult_202_n65, S => 
                           mult_202_n66);
   mult_202_U41 : ADFULD1 port map( A => mult_202_n92, B => mult_202_n98, CI =>
                           mult_202_n104, CO => mult_202_n63, S => mult_202_n64
                           );
   mult_202_U40 : ADFULD1 port map( A => mult_202_n67, B => mult_202_n111, CI 
                           => mult_202_n64, CO => mult_202_n61, S => 
                           mult_202_n62);
   mult_202_U39 : ADHALFDL port map( A => mult_202_n85, B => mult_202_n91, CO 
                           => mult_202_n59, S => mult_202_n60);
   mult_202_U38 : ADFULD1 port map( A => mult_202_n97, B => mult_202_n110, CI 
                           => mult_202_n103, CO => mult_202_n57, S => 
                           mult_202_n58);
   mult_202_U37 : ADFULD1 port map( A => mult_202_n63, B => mult_202_n60, CI =>
                           mult_202_n58, CO => mult_202_n55, S => mult_202_n56)
                           ;
   mult_202_U36 : ADHALFDL port map( A => mult_202_n96, B => mult_202_n90, CO 
                           => mult_202_n53, S => mult_202_n54);
   mult_202_U35 : ADFULD1 port map( A => mult_202_n84, B => mult_202_n102, CI 
                           => mult_202_n78, CO => mult_202_n51, S => 
                           mult_202_n52);
   mult_202_U34 : ADFULD1 port map( A => mult_202_n59, B => mult_202_n109, CI 
                           => mult_202_n54, CO => mult_202_n49, S => 
                           mult_202_n50);
   mult_202_U33 : ADFULD1 port map( A => mult_202_n52, B => mult_202_n57, CI =>
                           mult_202_n50, CO => mult_202_n47, S => mult_202_n48)
                           ;
   mult_202_U30 : ADFULD1 port map( A => mult_202_n101, B => mult_202_n89, CI 
                           => mult_202_n77, CO => mult_202_n43, S => 
                           mult_202_n44);
   mult_202_U29 : ADFULD1 port map( A => mult_202_n46, B => mult_202_n53, CI =>
                           mult_202_n51, CO => mult_202_n41, S => mult_202_n42)
                           ;
   mult_202_U28 : ADFULD1 port map( A => mult_202_n49, B => mult_202_n44, CI =>
                           mult_202_n42, CO => mult_202_n39, S => mult_202_n40)
                           ;
   mult_202_U26 : ADFULD1 port map( A => mult_202_n82, B => mult_202_n88, CI =>
                           mult_202_n76, CO => mult_202_n35, S => mult_202_n36)
                           ;
   mult_202_U25 : ADFULD1 port map( A => mult_202_n45, B => mult_202_n38, CI =>
                           mult_202_n43, CO => mult_202_n33, S => mult_202_n34)
                           ;
   mult_202_U24 : ADFULD1 port map( A => mult_202_n41, B => mult_202_n36, CI =>
                           mult_202_n34, CO => mult_202_n31, S => mult_202_n32)
                           ;
   mult_202_U23 : ADFULD1 port map( A => mult_202_n87, B => mult_202_n167, CI 
                           => mult_202_n75, CO => mult_202_n29, S => 
                           mult_202_n30);
   mult_202_U22 : ADFULD1 port map( A => mult_202_n94, B => mult_202_n81, CI =>
                           mult_202_n35, CO => mult_202_n27, S => mult_202_n28)
                           ;
   mult_202_U21 : ADFULD1 port map( A => mult_202_n33, B => mult_202_n30, CI =>
                           mult_202_n28, CO => mult_202_n25, S => mult_202_n26)
                           ;
   mult_202_U20 : ADFULD1 port map( A => mult_202_n86, B => mult_202_n80, CI =>
                           mult_202_n74, CO => mult_202_n23, S => mult_202_n24)
                           ;
   mult_202_U19 : ADFULD1 port map( A => mult_202_n24, B => mult_202_n29, CI =>
                           mult_202_n27, CO => mult_202_n21, S => mult_202_n22)
                           ;
   mult_202_U17 : ADFULD1 port map( A => mult_202_n20, B => mult_202_n73, CI =>
                           mult_202_n23, CO => mult_202_n17, S => mult_202_n18)
                           ;
   mult_202_U16 : ADFULD1 port map( A => mult_202_n79, B => mult_202_n168, CI 
                           => mult_202_n72, CO => mult_202_n15, S => 
                           mult_202_n16);
   mult_202_U15 : ADHALFDL port map( A => mult_202_n115, B => mult_202_n108, CO
                           => mult_202_n14, S => m_out_1_port);
   mult_202_U14 : ADFULD1 port map( A => mult_202_n114, B => mult_202_n107, CI 
                           => mult_202_n14, CO => mult_202_n13, S => 
                           m_out_2_port);
   mult_202_U13 : ADFULD1 port map( A => mult_202_n70, B => mult_202_n100, CI 
                           => mult_202_n13, CO => mult_202_n12, S => 
                           m_out_3_port);
   mult_202_U12 : ADFULD1 port map( A => mult_202_n66, B => mult_202_n68, CI =>
                           mult_202_n12, CO => mult_202_n11, S => m_out_4_port)
                           ;
   mult_202_U11 : ADFULD1 port map( A => mult_202_n62, B => mult_202_n65, CI =>
                           mult_202_n11, CO => mult_202_n10, S => m_out_5_port)
                           ;
   mult_202_U10 : ADFULD1 port map( A => mult_202_n56, B => mult_202_n61, CI =>
                           mult_202_n10, CO => mult_202_n9, S => m_out_6_port);
   mult_202_U9 : ADFULD1 port map( A => mult_202_n48, B => mult_202_n55, CI => 
                           mult_202_n9, CO => mult_202_n8, S => m_out_7_port);
   mult_202_U8 : ADFULD1 port map( A => mult_202_n40, B => mult_202_n47, CI => 
                           mult_202_n8, CO => mult_202_n7, S => m_out_8_port);
   mult_202_U7 : ADFULD1 port map( A => mult_202_n32, B => mult_202_n39, CI => 
                           mult_202_n7, CO => mult_202_n6, S => m_out_9_port);
   mult_202_U6 : ADFULD1 port map( A => mult_202_n26, B => mult_202_n31, CI => 
                           mult_202_n6, CO => mult_202_n5, S => m_out_10_port);
   mult_202_U5 : ADFULD1 port map( A => mult_202_n22, B => mult_202_n25, CI => 
                           mult_202_n5, CO => mult_202_n4, S => m_out_11_port);
   mult_202_U4 : ADFULD1 port map( A => mult_202_n21, B => mult_202_n18, CI => 
                           mult_202_n4, CO => mult_202_n3, S => m_out_12_port);
   mult_202_U3 : ADFULD1 port map( A => mult_202_n17, B => mult_202_n16, CI => 
                           mult_202_n3, CO => mult_202_n2, S => m_out_13_port);

end flat_rtl_none_10;
