
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_MAP1_overlapped is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type SIGNED is array (INTEGER range <>) of std_logic;

end CONV_PACK_MAP1_overlapped;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_MAP1_overlapped.all;

architecture hier_rtl_none_10 of MAP1_overlapped_DW_mult_tc_2 is

   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n29, n30, n31, n32, n33
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, product_6_port, product_7_port,
      product_8_port, product_9_port, product_10_port, product_11_port, 
      product_12_port, n119, product_13_port, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n_1003, n_1004, n_1005, n_1006, n_1007, 
      n_1008, n_1009, n_1010, n_1011 : std_logic;

begin
   product <= ( product_13_port, product_13_port, product_12_port, 
      product_11_port, product_10_port, product_9_port, product_8_port, 
      product_7_port, product_6_port, n_1003, n_1004, n_1005, n_1006, n_1007, 
      n_1008 );
   
   U4 : ADFULD1 port map( A => n12, B => n46, CI => n3, CO => n2, S => 
                           product_12_port);
   U5 : ADFULD1 port map( A => n13, B => n14, CI => n4, CO => n3, S => 
                           product_11_port);
   U6 : ADFULD1 port map( A => n15, B => n18, CI => n5, CO => n4, S => 
                           product_10_port);
   U7 : ADFULD1 port map( A => n19, B => n24, CI => n6, CO => n5, S => 
                           product_9_port);
   U8 : ADFULD1 port map( A => n25, B => n30, CI => n7, CO => n6, S => 
                           product_8_port);
   U9 : ADFULD1 port map( A => n31, B => n36, CI => n8, CO => n7, S => 
                           product_7_port);
   U10 : ADFULD1 port map( A => n37, B => n40, CI => n9, CO => n8, S => 
                           product_6_port);
   U11 : ADFULD1 port map( A => n10, B => n43, CI => n41, CO => n9, S => n_1009
                           );
   U12 : ADFULD1 port map( A => n11, B => n58, CI => n45, CO => n10, S => 
                           n_1010);
   U13 : ADHALFDL port map( A => n71, B => n66, CO => n11, S => n_1011);
   U14 : ADFULD1 port map( A => n51, B => n47, CI => n16, CO => n12, S => n13);
   U15 : ADFULD1 port map( A => n20, B => n48, CI => n17, CO => n14, S => n15);
   U16 : ADFULD1 port map( A => n52, B => n124, CI => n59, CO => n16, S => n17)
                           ;
   U17 : ADFULD1 port map( A => n26, B => n23, CI => n21, CO => n18, S => n19);
   U18 : ADFULD1 port map( A => n126, B => n60, CI => n53, CO => n20, S => n21)
                           ;
   U20 : ADFULD1 port map( A => n32, B => n29, CI => n27, CO => n24, S => n25);
   U21 : ADFULD1 port map( A => n128, B => n61, CI => n54, CO => n26, S => n27)
                           ;
   U23 : ADFULD1 port map( A => n38, B => n35, CI => n33, CO => n30, S => n31);
   U24 : ADFULD1 port map( A => n55, B => n62, CI => n67, CO => n32, S => n33);
   U26 : ADFULD1 port map( A => n42, B => n68, CI => n39, CO => n36, S => n37);
   U27 : ADFULD1 port map( A => n49, B => n56, CI => n63, CO => n38, S => n39);
   U28 : ADFULD1 port map( A => n64, B => n69, CI => n44, CO => n40, S => n41);
   U29 : ADHALFDL port map( A => n50, B => n57, CO => n42, S => n43);
   U30 : ADHALFDL port map( A => n65, B => n70, CO => n44, S => n45);
   U78 : INVD1 port map( A => a(3), Z => n119);
   U79 : INVD1 port map( A => n2, Z => product_13_port);
   U80 : INVD1 port map( A => b(4), Z => n123);
   U81 : INVD1 port map( A => b(2), Z => n127);
   U82 : INVD1 port map( A => b(3), Z => n125);
   U83 : INVD1 port map( A => n35, Z => n128);
   U84 : INVD1 port map( A => n29, Z => n126);
   U85 : INVD1 port map( A => n23, Z => n124);
   U86 : INVD1 port map( A => b(1), Z => n129);
   U87 : INVD1 port map( A => b(0), Z => n130);
   U88 : INVD1 port map( A => b(5), Z => n122);
   U89 : INVD1 port map( A => b(6), Z => n121);
   U90 : NOR2D1 port map( A1 => n119, A2 => n125, Z => n71);
   U91 : NOR2D1 port map( A1 => n119, A2 => n123, Z => n70);
   U92 : NOR2D1 port map( A1 => n119, A2 => n122, Z => n69);
   U93 : NOR2D1 port map( A1 => n119, A2 => n121, Z => n68);
   U94 : NAN2D1 port map( A1 => b(7), A2 => a(0), Z => n67);
   U95 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n66);
   U96 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n65);
   U97 : NOR2D1 port map( A1 => n127, A2 => n119, Z => n64);
   U98 : NOR2D1 port map( A1 => n125, A2 => n119, Z => n63);
   U99 : NOR2D1 port map( A1 => n123, A2 => n119, Z => n62);
   U100 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n61);
   U101 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n60);
   U102 : NAN2D1 port map( A1 => a(3), A2 => b(7), Z => n59);
   U103 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n58);
   U104 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n57);
   U105 : NOR2D1 port map( A1 => n127, A2 => n119, Z => n56);
   U106 : NOR2D1 port map( A1 => n125, A2 => n119, Z => n55);
   U107 : NOR2D1 port map( A1 => n123, A2 => n119, Z => n54);
   U108 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n53);
   U109 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n52);
   U110 : NAN2D1 port map( A1 => a(4), A2 => b(7), Z => n51);
   U111 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n50);
   U112 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n49);
   U113 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n48);
   U114 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n47);
   U115 : NAN2D1 port map( A1 => a(5), A2 => b(7), Z => n46);
   U116 : NAN2D1 port map( A1 => a(5), A2 => b(2), Z => n35);
   U117 : NAN2D1 port map( A1 => a(5), A2 => b(3), Z => n29);
   U118 : NAN2D1 port map( A1 => a(5), A2 => b(4), Z => n23);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_MAP1_overlapped.all;

architecture hier_rtl_none_10 of MAP1_overlapped_DW_mult_tc_1 is

   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n16, n17, n18, 
      n19, n20, n21, n23, n24, n25, n26, n27, n28, n29, n30, n32, n33, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n50, 
      n51, n52, n53, n54, n55, n56, n57, n60, n62, n63, n64, n65, n66, n67, n68
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, 
      n86, n87, n88, n89, n90, n91, n92, product_1_port, product_2_port, 
      product_3_port, product_4_port, product_5_port, product_6_port, 
      product_7_port, product_8_port, product_9_port, product_10_port, 
      product_11_port, product_12_port, product_13_port, product_14_port, n184,
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n_1014 : std_logic;

begin
   product <= ( n_1014, product_14_port, product_13_port, product_12_port, 
      product_11_port, product_10_port, product_9_port, product_8_port, 
      product_7_port, product_6_port, product_5_port, product_4_port, 
      product_3_port, product_2_port, product_1_port, b(0) );
   
   U3 : ADFULD1 port map( A => n17, B => n16, CI => n3, CO => n2, S => 
                           product_13_port);
   U4 : ADFULD1 port map( A => n19, B => n18, CI => n4, CO => n3, S => 
                           product_12_port);
   U5 : ADFULD1 port map( A => n20, B => n23, CI => n5, CO => n4, S => 
                           product_11_port);
   U6 : ADFULD1 port map( A => n24, B => n27, CI => n6, CO => n5, S => 
                           product_10_port);
   U7 : ADFULD1 port map( A => n28, B => n33, CI => n7, CO => n6, S => 
                           product_9_port);
   U8 : ADFULD1 port map( A => n34, B => n39, CI => n8, CO => n7, S => 
                           product_8_port);
   U9 : ADFULD1 port map( A => n40, B => n45, CI => n9, CO => n8, S => 
                           product_7_port);
   U10 : ADFULD1 port map( A => n46, B => n185, CI => n10, CO => n9, S => 
                           product_6_port);
   U11 : ADFULD1 port map( A => n50, B => n52, CI => n11, CO => n10, S => 
                           product_5_port);
   U12 : ADFULD1 port map( A => n54, B => n55, CI => n12, CO => n11, S => 
                           product_4_port);
   U13 : ADFULD1 port map( A => n56, B => n83, CI => n184, CO => n12, S => 
                           product_3_port);
   U15 : ADHALFDL port map( A => n92, B => n60, CO => n14, S => product_1_port)
                           ;
   U17 : ADFULD1 port map( A => n62, B => n21, CI => n69, CO => n17, S => n18);
   U18 : ADFULD1 port map( A => n190, B => n63, CI => n25, CO => n19, S => n20)
                           ;
   U20 : ADFULD1 port map( A => n29, B => n77, CI => n26, CO => n23, S => n24);
   U21 : ADFULD1 port map( A => n70, B => n191, CI => n64, CO => n25, S => n26)
                           ;
   U22 : ADFULD1 port map( A => n35, B => n37, CI => n30, CO => n27, S => n28);
   U23 : ADFULD1 port map( A => n65, B => n71, CI => n32, CO => n29, S => n30);
   U25 : ADFULD1 port map( A => n41, B => n38, CI => n36, CO => n33, S => n34);
   U26 : ADFULD1 port map( A => n66, B => n72, CI => n43, CO => n35, S => n36);
   U29 : ADFULD1 port map( A => n44, B => n47, CI => n42, CO => n39, S => n40);
   U30 : ADFULD1 port map( A => n67, B => n73, CI => n57, CO => n41, S => n42);
   U31 : ADHALFDL port map( A => n79, B => n86, CO => n43, S => n44);
   U32 : ADFULD1 port map( A => n51, B => n74, CI => n48, CO => n45, S => n46);
   U33 : ADFULD1 port map( A => n68, B => n87, CI => n80, CO => n47, S => n48);
   U35 : ADHALFDL port map( A => n81, B => n88, CO => n51, S => n52);
   U36 : ADFULD1 port map( A => n89, B => n76, CI => n82, CO => n53, S => n54);
   U37 : ADHALFDL port map( A => n186, B => n90, CO => n55, S => n56);
   U135 : AND2D1 port map( A1 => n14, A2 => n91, Z => n184);
   U136 : INVD1 port map( A => n205, Z => n195);
   U137 : AND2D1 port map( A1 => n53, A2 => n75, Z => n185);
   U138 : INVD1 port map( A => a(6), Z => n186);
   U139 : EXOR2D1 port map( A1 => a(6), A2 => n187, Z => n205);
   U140 : INVD1 port map( A => a(4), Z => n187);
   U141 : NAN2D1 port map( A1 => n193, A2 => n186, Z => n212);
   U142 : NAN2D1 port map( A1 => n192, A2 => n186, Z => n32);
   U143 : NAN2D1 port map( A1 => n186, A2 => n188, Z => n77);
   U144 : NOR2D1 port map( A1 => a(5), A2 => n203, Z => n70);
   U145 : INVD1 port map( A => n32, Z => n191);
   U146 : NOR2D1 port map( A1 => n205, A2 => n209, Z => n64);
   U147 : NOR2D1 port map( A1 => a(5), A2 => n204, Z => n21);
   U148 : NAN2D1 port map( A1 => n187, A2 => n189, Z => n69);
   U149 : NOR2D1 port map( A1 => n205, A2 => n211, Z => n62);
   U150 : INVD1 port map( A => n204, Z => n189);
   U151 : NAN2D1 port map( A1 => n195, A2 => n197, Z => n16);
   U152 : NAN2D1 port map( A1 => n195, A2 => n197, Z => n196);
   U153 : NOR2D1 port map( A1 => b(0), A2 => a(6), Z => n83);
   U154 : NOR2D1 port map( A1 => a(5), A2 => n199, Z => n74);
   U155 : NOR2D1 port map( A1 => b(3), A2 => a(6), Z => n80);
   U156 : NOR2D1 port map( A1 => b(1), A2 => a(6), Z => n82);
   U157 : NOR2D1 port map( A1 => a(5), A2 => n200, Z => n73);
   U158 : NOR3D1 port map( A1 => n205, A2 => n186, A3 => b(0), Z => n57);
   U159 : NOR2D1 port map( A1 => n205, A2 => n206, Z => n67);
   U160 : NOR2D1 port map( A1 => b(2), A2 => a(6), Z => n81);
   U161 : NOR2D1 port map( A1 => a(5), A2 => n198, Z => n75);
   U162 : NOR2D1 port map( A1 => b(4), A2 => a(6), Z => n79);
   U163 : NOR2D1 port map( A1 => a(5), A2 => n201, Z => n72);
   U164 : NOR2D1 port map( A1 => n205, A2 => n207, Z => n66);
   U165 : NOR2D1 port map( A1 => a(5), A2 => n202, Z => n71);
   U166 : NOR2D1 port map( A1 => n205, A2 => n208, Z => n65);
   U167 : INVD1 port map( A => b(0), Z => n194);
   U168 : INVD1 port map( A => b(6), Z => n192);
   U169 : INVD1 port map( A => b(5), Z => n193);
   U170 : INVD1 port map( A => n21, Z => n190);
   U171 : NOR2D1 port map( A1 => n205, A2 => n210, Z => n63);
   U172 : INVD1 port map( A => b(7), Z => n188);
   U173 : EXOR2D1 port map( A1 => n75, A2 => n53, Z => n50);
   U174 : EXOR2D1 port map( A1 => n91, A2 => n14, Z => product_2_port);
   U175 : EXNOR3D1 port map( A1 => n2, A2 => n16, A3 => n196, Z => 
                           product_14_port);
   U176 : EXOR2D1 port map( A1 => b(1), A2 => a(1), Z => n92);
   U177 : EXOR2D1 port map( A1 => b(2), A2 => a(1), Z => n91);
   U178 : EXOR2D1 port map( A1 => b(3), A2 => a(1), Z => n90);
   U179 : EXOR2D1 port map( A1 => b(4), A2 => a(1), Z => n89);
   U180 : EXNOR2D1 port map( A1 => n193, A2 => a(1), Z => n88);
   U181 : EXNOR2D1 port map( A1 => n192, A2 => a(1), Z => n87);
   U182 : NOR2D1 port map( A1 => a(5), A2 => n194, Z => n76);
   U183 : EXNOR2D1 port map( A1 => b(1), A2 => a(5), Z => n198);
   U184 : EXNOR2D1 port map( A1 => b(2), A2 => a(5), Z => n199);
   U185 : EXNOR2D1 port map( A1 => b(3), A2 => a(5), Z => n200);
   U186 : EXNOR2D1 port map( A1 => b(4), A2 => a(5), Z => n201);
   U187 : EXNOR2D1 port map( A1 => b(5), A2 => a(5), Z => n202);
   U188 : NOR2D1 port map( A1 => n205, A2 => n194, Z => n68);
   U189 : EXNOR2D1 port map( A1 => b(1), A2 => a(7), Z => n206);
   U190 : EXNOR2D1 port map( A1 => b(2), A2 => a(7), Z => n207);
   U191 : EXNOR2D1 port map( A1 => b(3), A2 => a(7), Z => n208);
   U192 : EXNOR2D1 port map( A1 => b(4), A2 => a(7), Z => n209);
   U193 : EXNOR2D1 port map( A1 => b(5), A2 => a(7), Z => n210);
   U194 : NOR2M1D1 port map( A1 => a(1), A2 => b(0), Z => n60);
   U195 : EXNOR2D1 port map( A1 => n212, A2 => n86, Z => n38);
   U196 : NAN2D1 port map( A1 => n212, A2 => n86, Z => n37);
   U197 : EXNOR2D1 port map( A1 => n188, A2 => a(1), Z => n86);
   U198 : EXOR2D1 port map( A1 => b(6), A2 => n187, Z => n203);
   U199 : EXNOR2D1 port map( A1 => b(7), A2 => a(5), Z => n204);
   U200 : EXOR2D1 port map( A1 => b(6), A2 => n186, Z => n211);
   U201 : EXNOR2D1 port map( A1 => b(7), A2 => n186, Z => n197);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_MAP1_overlapped.all;

architecture hier_rtl_none_10 of MAP1_overlapped_DW_mult_tc_0 is

   component MUX2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIEHI
      port( Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n18, n19, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n34, n35
      , n36, n37, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n126, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n185, n186, n187 : std_logic;

begin
   
   U3 : ADFULD1 port map( A => n18, B => n175, CI => n3, CO => n2, S => 
                           product(13));
   U4 : ADFULD1 port map( A => n20, B => n19, CI => n4, CO => n3, S => 
                           product(12));
   U5 : ADFULD1 port map( A => n21, B => n24, CI => n5, CO => n4, S => 
                           product(11));
   U6 : ADFULD1 port map( A => n25, B => n28, CI => n6, CO => n5, S => 
                           product(10));
   U7 : ADFULD1 port map( A => n29, B => n34, CI => n7, CO => n6, S => 
                           product(9));
   U8 : ADFULD1 port map( A => n35, B => n39, CI => n8, CO => n7, S => 
                           product(8));
   U9 : ADFULD1 port map( A => n40, B => n43, CI => n9, CO => n8, S => 
                           product(7));
   U10 : ADFULD1 port map( A => n44, B => n47, CI => n10, CO => n9, S => 
                           product(6));
   U11 : ADFULD1 port map( A => n48, B => n49, CI => n11, CO => n10, S => 
                           product(5));
   U12 : ADFULD1 port map( A => n50, B => n51, CI => n12, CO => n11, S => 
                           product(4));
   U13 : ADFULD1 port map( A => n52, B => n53, CI => n13, CO => n12, S => 
                           product(3));
   U14 : ADFULD1 port map( A => n14, B => n105, CI => n54, CO => n13, S => 
                           product(2));
   U15 : ADHALFDL port map( A => n112, B => n15, CO => n14, S => product(1));
   U18 : ADFULD1 port map( A => n82, B => n88, CI => n22, CO => n18, S => n19);
   U19 : ADFULD1 port map( A => n178, B => n89, CI => n26, CO => n20, S => n21)
                           ;
   U21 : ADFULD1 port map( A => n30, B => n90, CI => n27, CO => n24, S => n25);
   U22 : ADFULD1 port map( A => n97, B => b(7), CI => n83, CO => n26, S => n27)
                           ;
   U23 : ADFULD1 port map( A => n36, B => n91, CI => n31, CO => n28, S => n29);
   U24 : ADFULD1 port map( A => n98, B => n176, CI => n84, CO => n30, S => n31)
                           ;
   U26 : ADFULD1 port map( A => n41, B => n92, CI => n37, CO => n34, S => n35);
   U27 : ADFULD1 port map( A => n99, B => n176, CI => n85, CO => n36, S => n37)
                           ;
   U29 : ADFULD1 port map( A => n45, B => n93, CI => n42, CO => n39, S => n40);
   U30 : ADFULD1 port map( A => n100, B => n106, CI => n86, CO => n41, S => n42
                           );
   U31 : ADFULD1 port map( A => n94, B => n87, CI => n46, CO => n43, S => n44);
   U32 : ADFULD1 port map( A => a(7), B => n107, CI => n101, CO => n45, S => 
                           n46);
   U33 : ADFULD1 port map( A => n102, B => n108, CI => n95, CO => n47, S => n48
                           );
   U34 : ADFULD1 port map( A => n103, B => n109, CI => n96, CO => n49, S => n50
                           );
   U35 : ADHALFDL port map( A => n104, B => n110, CO => n51, S => n52);
   U36 : ADHALFDL port map( A => n111, B => a(3), CO => n53, S => n54);
   U39 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n55, Z => n16);
   U41 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n56, Z => n82);
   U43 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n57, Z => n22);
   U45 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n58, Z => n83);
   U47 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n59, Z => n84);
   U49 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n60, Z => n85);
   U51 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n61, Z => n86);
   U53 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n62, Z => n87);
   U56 : NOR2D1 port map( A1 => n177, A2 => n174, Z => n89);
   U58 : NOR2D1 port map( A1 => n179, A2 => n174, Z => n90);
   U60 : NOR2D1 port map( A1 => n180, A2 => n174, Z => n91);
   U62 : NOR2D1 port map( A1 => n181, A2 => n174, Z => n92);
   U64 : NOR2D1 port map( A1 => n182, A2 => n174, Z => n93);
   U66 : NOR2D1 port map( A1 => n183, A2 => n174, Z => n94);
   U68 : NOR2D1 port map( A1 => n185, A2 => n174, Z => n95);
   U70 : NOR2D1 port map( A1 => n186, A2 => n174, Z => n96);
   U74 : EXNOR2D1 port map( A1 => a(3), A2 => n176, Z => n98);
   U76 : EXNOR2D1 port map( A1 => a(3), A2 => n177, Z => n99);
   U78 : EXNOR2D1 port map( A1 => a(3), A2 => n179, Z => n100);
   U80 : EXNOR2D1 port map( A1 => a(3), A2 => n180, Z => n101);
   U82 : EXNOR2D1 port map( A1 => a(3), A2 => n181, Z => n102);
   U84 : EXNOR2D1 port map( A1 => a(3), A2 => n182, Z => n103);
   U86 : EXNOR2D1 port map( A1 => a(3), A2 => n183, Z => n104);
   U88 : EXNOR2D1 port map( A1 => a(3), A2 => n185, Z => n105);
   U126 : INVD1 port map( A => a(7), Z => n174);
   U127 : NAN2D1 port map( A1 => a(6), A2 => n174, Z => n126);
   U128 : INVD1 port map( A => n16, Z => n175);
   U129 : INVD1 port map( A => n22, Z => n178);
   U130 : INVD1 port map( A => n15, Z => product(0));
   U131 : INVD1 port map( A => b(0), Z => n185);
   U132 : INVD1 port map( A => b(1), Z => n183);
   U133 : INVD1 port map( A => b(2), Z => n182);
   U134 : INVD1 port map( A => b(3), Z => n181);
   U135 : INVD1 port map( A => b(4), Z => n180);
   U136 : INVD1 port map( A => b(5), Z => n179);
   U137 : INVD1 port map( A => b(6), Z => n177);
   U138 : INVD1 port map( A => b(7), Z => n176);
   U139 : TIEHI port map( Z => n186);
   U140 : EXNOR3D1 port map( A1 => n2, A2 => n16, A3 => n187, Z => product(14))
                           ;
   U141 : MUXB2DL port map( A0 => n126, A1 => n174, SL => n176, Z => n187);
   U142 : EXNOR2D1 port map( A1 => a(3), A2 => b(7), Z => n97);
   U143 : NAN2M1D1 port map( A1 => n174, A2 => b(7), Z => n88);
   U144 : NAN2D1 port map( A1 => a(6), A2 => b(0), Z => n62);
   U145 : MUX2DL port map( A0 => n185, A1 => n183, SL => a(6), Z => n61);
   U146 : MUX2DL port map( A0 => n183, A1 => n182, SL => a(6), Z => n60);
   U147 : MUX2DL port map( A0 => n182, A1 => n181, SL => a(6), Z => n59);
   U148 : MUX2DL port map( A0 => n181, A1 => n180, SL => a(6), Z => n58);
   U149 : MUX2DL port map( A0 => n180, A1 => n179, SL => a(6), Z => n57);
   U150 : MUX2DL port map( A0 => n179, A1 => n177, SL => a(6), Z => n56);
   U151 : MUX2DL port map( A0 => n177, A1 => n176, SL => a(6), Z => n55);
   U152 : NAN2D1 port map( A1 => a(0), A2 => b(0), Z => n15);
   U153 : MUX2DL port map( A0 => n185, A1 => n183, SL => a(0), Z => n112);
   U154 : MUX2DL port map( A0 => n183, A1 => n182, SL => a(0), Z => n111);
   U155 : MUX2DL port map( A0 => n182, A1 => n181, SL => a(0), Z => n110);
   U156 : MUX2DL port map( A0 => n181, A1 => n180, SL => a(0), Z => n109);
   U157 : MUX2DL port map( A0 => n180, A1 => n179, SL => a(0), Z => n108);
   U158 : MUX2DL port map( A0 => n179, A1 => n177, SL => a(0), Z => n107);
   U159 : MUX2DL port map( A0 => n177, A1 => n176, SL => a(0), Z => n106);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_MAP1_overlapped.all;

architecture hier_rtl_none_10 of MAP1_overlapped_DW01_add_3 is

   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, n1
      , n2, n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1_13 : ADFULD1 port map( A => A(13), B => B(13), CI => carry_13_port, CO =>
                           carry_14_port, S => SUM(13));
   U1_12 : ADFULD1 port map( A => A(12), B => B(12), CI => carry_12_port, CO =>
                           carry_13_port, S => SUM(12));
   U1_11 : ADFULD1 port map( A => A(11), B => B(11), CI => carry_11_port, CO =>
                           carry_12_port, S => SUM(11));
   U1_10 : ADFULD1 port map( A => A(10), B => B(10), CI => carry_10_port, CO =>
                           carry_11_port, S => SUM(10));
   U1_9 : ADFULD1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : ADFULD1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : ADFULD1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : ADFULD1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_14 : EXOR3D1 port map( A1 => A(14), A2 => B(14), A3 => carry_14_port, Z 
                           => SUM(14));
   U1 : OAI21M20D1 port map( A1 => n1, A2 => A(5), B => n2, Z => carry_6_port);
   U2 : OAI21D1 port map( A1 => A(5), A2 => n1, B => B(5), Z => n2);
   U3 : OAI21M20D1 port map( A1 => n3, A2 => A(4), B => n4, Z => n1);
   U4 : OAI21D1 port map( A1 => A(4), A2 => n3, B => B(4), Z => n4);
   U5 : OAI21M20D1 port map( A1 => n5, A2 => A(3), B => n6, Z => n3);
   U6 : OAI21D1 port map( A1 => A(3), A2 => n5, B => B(3), Z => n6);
   U7 : OAI21M20D1 port map( A1 => n7, A2 => A(2), B => n8, Z => n5);
   U8 : OAI21D1 port map( A1 => A(2), A2 => n7, B => B(2), Z => n8);
   U9 : OAI21M20D1 port map( A1 => A(1), A2 => B(1), B => n9, Z => n7);
   U10 : OAI211D1 port map( A1 => A(1), A2 => B(1), B => A(0), C => B(0), Z => 
                           n9);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_MAP1_overlapped.all;

architecture hier_rtl_none_10 of MAP1_overlapped is

   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIEHI
      port( Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component MAP1_overlapped_DW_mult_tc_0
      port( a, b : in std_logic_vector (7 downto 0);  product : out 
            std_logic_vector (15 downto 0));
   end component;
   
   component MAP1_overlapped_DW_mult_tc_1
      port( a, b : in std_logic_vector (7 downto 0);  product : out 
            std_logic_vector (15 downto 0));
   end component;
   
   component MAP1_overlapped_DW_mult_tc_2
      port( a : in std_logic_vector (6 downto 0);  b : in std_logic_vector (7 
            downto 0);  product : out std_logic_vector (14 downto 0));
   end component;
   
   component MAP1_overlapped_DW01_add_3
      port( A, B : in std_logic_vector (14 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (14 downto 0);  CO : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal arx_i1_reg_7_port, arx_i1_reg_6_port, arx_i1_reg_5_port, 
      arx_i1_reg_4_port, arx_i1_reg_3_port, arx_i1_reg_2_port, 
      arx_i1_reg_1_port, arx_i1_reg_0_port, arx_r1_reg_14_port, 
      arx_r1_reg_13_port, arx_r1_reg_12_port, arx_r1_reg_11_port, 
      arx_r1_reg_10_port, arx_r1_reg_9_port, arx_r1_reg_8_port, 
      arx_r1_reg_7_port, arx_r1_reg_6_port, arx_r1_reg_5_port, 
      arx_r1_reg_4_port, arx_r1_reg_3_port, arx_r1_reg_2_port, 
      arx_r1_reg_1_port, arx_r1_reg_0_port, arx_r2_reg_14_port, 
      arx_r2_reg_13_port, arx_r2_reg_12_port, arx_r2_reg_11_port, 
      arx_r2_reg_10_port, arx_r2_reg_9_port, arx_r2_reg_8_port, 
      arx_r2_reg_7_port, arx_r2_reg_6_port, arx_r2_reg_5_port, 
      arx_r2_reg_4_port, arx_r2_reg_3_port, arx_r2_reg_2_port, 
      arx_r2_reg_1_port, arx_r2_reg_0_port, arx_r3_reg_14_port, 
      arx_r3_reg_13_port, arx_r3_reg_12_port, arx_r3_reg_11_port, 
      arx_r3_reg_10_port, arx_r3_reg_9_port, arx_r3_reg_8_port, 
      arx_r3_reg_7_port, arx_r4_reg_14_port, arx_r4_reg_13_port, 
      arx_r4_reg_12_port, arx_r4_reg_11_port, arx_r4_reg_10_port, 
      arx_r4_reg_9_port, arx_r4_reg_8_port, arx_r4_reg_7_port, 
      arx_r4_reg_6_port, arx_state_reg_1_port, arx_state_reg_0_port, 
      m1_in_r_7_port, m1_in_r_6_port, m1_in_r_5_port, m1_in_r_4_port, 
      m1_in_r_3_port, m1_in_r_2_port, m1_in_r_1_port, m1_in_r_0_port, 
      m1_out_14_port, m1_out_13_port, m1_out_12_port, m1_out_11_port, 
      m1_out_10_port, m1_out_9_port, m1_out_8_port, m1_out_7_port, 
      m1_out_6_port, m1_out_5_port, m1_out_4_port, m1_out_3_port, m1_out_2_port
      , m1_out_1_port, m1_out_0_port, m2_in_l_5_port, m2_in_r_7_port, 
      m2_in_r_6_port, m2_in_r_5_port, m2_in_r_4_port, m2_in_r_3_port, 
      m2_in_r_2_port, m2_in_r_1_port, m2_in_r_0_port, m2_out_14_port, 
      m2_out_13_port, m2_out_12_port, m2_out_11_port, m2_out_10_port, 
      m2_out_9_port, m2_out_8_port, m2_out_7_port, m2_out_6_port, m2_out_5_port
      , m2_out_4_port, m2_out_3_port, m2_out_2_port, m2_out_1_port, 
      m2_out_0_port, m3_in_l_0, m3_in_r_7_port, m3_in_r_6_port, m3_in_r_5_port,
      m3_in_r_4_port, m3_in_r_3_port, m3_in_r_2_port, m3_in_r_1_port, 
      m3_in_r_0_port, m3_out_15, m3_out_13_port, m3_out_12_port, m3_out_11_port
      , m3_out_10_port, m3_out_9_port, m3_out_8_port, m3_out_7_port, 
      m3_out_6_port, a1_in_l_14_port, a1_in_l_13_port, a1_in_l_12_port, 
      a1_in_l_11_port, a1_in_l_10_port, a1_in_l_9_port, a1_in_l_8_port, 
      a1_in_l_7_port, a1_in_r_14_port, a1_in_r_13_port, a1_in_r_12_port, 
      a1_in_r_11_port, a1_in_r_10_port, a1_in_r_9_port, a1_in_r_8_port, 
      a1_in_r_7_port, a1_in_r_6_port, a1_in_r_5_port, a1_in_r_4_port, 
      a1_in_r_3_port, a1_in_r_2_port, a1_in_r_1_port, a1_in_r_0_port, 
      a1_out_7_port, a1_out_6_port, a1_out_5_port, a1_out_4_port, a1_out_3_port
      , a1_out_2_port, a1_out_1_port, a1_out_0_port, a2_in_l_14_port, 
      a2_in_l_13_port, a2_in_l_12_port, a2_in_l_11_port, a2_in_l_10_port, 
      a2_in_l_9_port, a2_in_l_8_port, a2_in_l_7_port, a2_in_r_14_port, 
      a2_in_r_13_port, a2_in_r_12_port, a2_in_r_11_port, a2_in_r_10_port, 
      a2_in_r_9_port, a2_in_r_8_port, a2_in_r_7_port, a2_out_7_port, 
      a2_out_6_port, a2_out_5_port, a2_out_4_port, a2_out_3_port, a2_out_2_port
      , a2_out_1_port, a2_out_0_port, state_1_port, N106, N107, N108, N109, 
      N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, 
      N122, N123, N137, n55, n56, n57, n58, n60, n61, n62, n63, n64, n65, n66, 
      n67, n68, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n91, n92, add_416_C224_rn_carry_1_port, add_416_C224_rn_carry_2_port, 
      add_416_C224_rn_carry_3_port, add_416_C224_rn_carry_4_port, 
      add_416_C224_rn_carry_5_port, add_416_C224_rn_carry_6_port, 
      add_416_C224_rn_carry_7_port, add_224_carry_8_port, add_224_carry_9_port,
      add_224_carry_10_port, add_224_carry_11_port, add_224_carry_12_port, 
      add_224_carry_13_port, add_224_carry_14_port, 
      add_416_C223_rn_carry_1_port, add_416_C223_rn_carry_2_port, 
      add_416_C223_rn_carry_3_port, add_416_C223_rn_carry_4_port, 
      add_416_C223_rn_carry_5_port, add_416_C223_rn_carry_6_port, 
      add_416_C223_rn_carry_7_port, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n1060, n1070, n1080, n1090, n1100, n1110, 
      n1120, n1130, n1140, n1150, n1160, n1170, n1180, n1190, n_1027, n_1028, 
      n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, 
      n_1038, n_1039, n_1040, n_1041 : std_logic;

begin
   
   U119 : OAI21D1 port map( A1 => n1060, A2 => n1170, B => n58, Z => n78);
   U120 : AOI22D1 port map( A1 => n104, A2 => a1_out_7_port, B1 => 
                           m2_out_14_port, B2 => n60, Z => n58);
   U121 : OAI21D1 port map( A1 => n1060, A2 => n1160, B => n61, Z => n79);
   U122 : AOI22D1 port map( A1 => n104, A2 => a1_out_6_port, B1 => 
                           m2_out_13_port, B2 => n60, Z => n61);
   U123 : OAI21D1 port map( A1 => n1060, A2 => n1150, B => n62, Z => n80);
   U124 : AOI22D1 port map( A1 => n104, A2 => a1_out_5_port, B1 => 
                           m2_out_12_port, B2 => n60, Z => n62);
   U125 : OAI21D1 port map( A1 => n1060, A2 => n1140, B => n63, Z => n81);
   U126 : AOI22D1 port map( A1 => n104, A2 => a1_out_4_port, B1 => 
                           m2_out_11_port, B2 => n60, Z => n63);
   U127 : OAI21D1 port map( A1 => n1060, A2 => n1130, B => n64, Z => n82);
   U128 : AOI22D1 port map( A1 => n104, A2 => a1_out_3_port, B1 => 
                           m2_out_10_port, B2 => n60, Z => n64);
   U129 : OAI21D1 port map( A1 => n1060, A2 => n1120, B => n65, Z => n83);
   U130 : AOI22D1 port map( A1 => n104, A2 => a1_out_2_port, B1 => 
                           m2_out_9_port, B2 => n60, Z => n65);
   U131 : OAI21D1 port map( A1 => n1060, A2 => n1110, B => n66, Z => n84);
   U132 : AOI22D1 port map( A1 => n104, A2 => a1_out_1_port, B1 => 
                           m2_out_8_port, B2 => n60, Z => n66);
   U133 : OAI21D1 port map( A1 => n1060, A2 => n1100, B => n67, Z => n85);
   U134 : AOI22D1 port map( A1 => n104, A2 => a1_out_0_port, B1 => 
                           m2_out_7_port, B2 => n60, Z => n67);
   add_223 : MAP1_overlapped_DW01_add_3 port map( A(14) => a1_in_l_14_port, 
                           A(13) => a1_in_l_13_port, A(12) => a1_in_l_12_port, 
                           A(11) => a1_in_l_11_port, A(10) => a1_in_l_10_port, 
                           A(9) => a1_in_l_9_port, A(8) => a1_in_l_8_port, A(7)
                           => a1_in_l_7_port, A(6) => n98, A(5) => n101, A(4) 
                           => n97, A(3) => n96, A(2) => n95, A(1) => n93, A(0) 
                           => n94, B(14) => a1_in_r_14_port, B(13) => 
                           a1_in_r_13_port, B(12) => a1_in_r_12_port, B(11) => 
                           a1_in_r_11_port, B(10) => a1_in_r_10_port, B(9) => 
                           a1_in_r_9_port, B(8) => a1_in_r_8_port, B(7) => 
                           a1_in_r_7_port, B(6) => a1_in_r_6_port, B(5) => 
                           a1_in_r_5_port, B(4) => a1_in_r_4_port, B(3) => 
                           a1_in_r_3_port, B(2) => a1_in_r_2_port, B(1) => 
                           a1_in_r_1_port, B(0) => a1_in_r_0_port, CI => n1190,
                           SUM(14) => N114, SUM(13) => N113, SUM(12) => N112, 
                           SUM(11) => N111, SUM(10) => N110, SUM(9) => N109, 
                           SUM(8) => N108, SUM(7) => N107, SUM(6) => N106, 
                           SUM(5) => n_1027, SUM(4) => n_1028, SUM(3) => n_1029
                           , SUM(2) => n_1030, SUM(1) => n_1031, SUM(0) => 
                           n_1032, CO => n_1033);
   mult_222 : MAP1_overlapped_DW_mult_tc_2 port map( a(6) => n1190, a(5) => 
                           m3_in_l_0, a(4) => m3_in_l_0, a(3) => m3_in_l_0, 
                           a(2) => n1190, a(1) => n1190, a(0) => m3_in_l_0, 
                           b(7) => m3_in_r_7_port, b(6) => m3_in_r_6_port, b(5)
                           => m3_in_r_5_port, b(4) => m3_in_r_4_port, b(3) => 
                           m3_in_r_3_port, b(2) => m3_in_r_2_port, b(1) => 
                           m3_in_r_1_port, b(0) => m3_in_r_0_port, product(14) 
                           => m3_out_15, product(13) => m3_out_13_port, 
                           product(12) => m3_out_12_port, product(11) => 
                           m3_out_11_port, product(10) => m3_out_10_port, 
                           product(9) => m3_out_9_port, product(8) => 
                           m3_out_8_port, product(7) => m3_out_7_port, 
                           product(6) => m3_out_6_port, product(5) => n_1034, 
                           product(4) => n_1035, product(3) => n_1036, 
                           product(2) => n_1037, product(1) => n_1038, 
                           product(0) => n_1039);
   mult_221 : MAP1_overlapped_DW_mult_tc_1 port map( a(7) => m3_in_l_0, a(6) =>
                           m3_in_l_0, a(5) => m2_in_l_5_port, a(4) => 
                           m2_in_l_5_port, a(3) => n1180, a(2) => m3_in_l_0, 
                           a(1) => m3_in_l_0, a(0) => n1180, b(7) => 
                           m2_in_r_7_port, b(6) => m2_in_r_6_port, b(5) => 
                           m2_in_r_5_port, b(4) => m2_in_r_4_port, b(3) => 
                           m2_in_r_3_port, b(2) => m2_in_r_2_port, b(1) => 
                           m2_in_r_1_port, b(0) => m2_in_r_0_port, product(15) 
                           => n_1040, product(14) => m2_out_14_port, 
                           product(13) => m2_out_13_port, product(12) => 
                           m2_out_12_port, product(11) => m2_out_11_port, 
                           product(10) => m2_out_10_port, product(9) => 
                           m2_out_9_port, product(8) => m2_out_8_port, 
                           product(7) => m2_out_7_port, product(6) => 
                           m2_out_6_port, product(5) => m2_out_5_port, 
                           product(4) => m2_out_4_port, product(3) => 
                           m2_out_3_port, product(2) => m2_out_2_port, 
                           product(1) => m2_out_1_port, product(0) => 
                           m2_out_0_port);
   mult_220 : MAP1_overlapped_DW_mult_tc_0 port map( a(7) => m2_in_l_5_port, 
                           a(6) => m3_in_l_0, a(5) => n1190, a(4) => 
                           m2_in_l_5_port, a(3) => m2_in_l_5_port, a(2) => 
                           n1190, a(1) => n1180, a(0) => m3_in_l_0, b(7) => 
                           m1_in_r_7_port, b(6) => m1_in_r_6_port, b(5) => 
                           m1_in_r_5_port, b(4) => m1_in_r_4_port, b(3) => 
                           m1_in_r_3_port, b(2) => m1_in_r_2_port, b(1) => 
                           m1_in_r_1_port, b(0) => m1_in_r_0_port, product(15) 
                           => n_1041, product(14) => m1_out_14_port, 
                           product(13) => m1_out_13_port, product(12) => 
                           m1_out_12_port, product(11) => m1_out_11_port, 
                           product(10) => m1_out_10_port, product(9) => 
                           m1_out_9_port, product(8) => m1_out_8_port, 
                           product(7) => m1_out_7_port, product(6) => 
                           m1_out_6_port, product(5) => m1_out_5_port, 
                           product(4) => m1_out_4_port, product(3) => 
                           m1_out_3_port, product(2) => m1_out_2_port, 
                           product(1) => m1_out_1_port, product(0) => 
                           m1_out_0_port);
   add_224_U1_8 : ADFULD1 port map( A => a2_in_l_8_port, B => a2_in_r_8_port, 
                           CI => add_224_carry_8_port, CO => 
                           add_224_carry_9_port, S => N117);
   add_224_U1_9 : ADFULD1 port map( A => a2_in_l_9_port, B => a2_in_r_9_port, 
                           CI => add_224_carry_9_port, CO => 
                           add_224_carry_10_port, S => N118);
   add_224_U1_10 : ADFULD1 port map( A => a2_in_l_10_port, B => a2_in_r_10_port
                           , CI => add_224_carry_10_port, CO => 
                           add_224_carry_11_port, S => N119);
   add_224_U1_11 : ADFULD1 port map( A => a2_in_l_11_port, B => a2_in_r_11_port
                           , CI => add_224_carry_11_port, CO => 
                           add_224_carry_12_port, S => N120);
   add_224_U1_12 : ADFULD1 port map( A => a2_in_l_12_port, B => a2_in_r_12_port
                           , CI => add_224_carry_12_port, CO => 
                           add_224_carry_13_port, S => N121);
   add_224_U1_13 : ADFULD1 port map( A => a2_in_l_13_port, B => a2_in_r_13_port
                           , CI => add_224_carry_13_port, CO => 
                           add_224_carry_14_port, S => N122);
   arx_r3_reg_reg_14_inst : DFERPQ1 port map( D => a1_out_7_port, CEB => n1060,
                           CK => clock, RB => resetn, Q => arx_r3_reg_14_port);
   arx_r4_reg_reg_14_inst : DFERPQ1 port map( D => m3_out_15, CEB => n1070, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_14_port);
   arx_r2_reg_reg_14_inst : DFFRPQ1 port map( D => n78, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_14_port);
   arx_r1_reg_reg_14_inst : DFERPQ1 port map( D => m1_out_14_port, CEB => n105,
                           CK => clock, RB => resetn, Q => arx_r1_reg_14_port);
   arx_i1_reg_reg_7_inst : DFERPQ1 port map( D => data_in(7), CEB => n56, CK =>
                           clock, RB => resetn, Q => arx_i1_reg_7_port);
   arx_r3_reg_reg_13_inst : DFERPQ1 port map( D => a1_out_6_port, CEB => n1060,
                           CK => clock, RB => resetn, Q => arx_r3_reg_13_port);
   arx_r4_reg_reg_13_inst : DFERPQ1 port map( D => m3_out_13_port, CEB => n1070
                           , CK => clock, RB => resetn, Q => arx_r4_reg_13_port
                           );
   arx_r2_reg_reg_13_inst : DFFRPQ1 port map( D => n79, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_13_port);
   arx_r1_reg_reg_13_inst : DFERPQ1 port map( D => m1_out_13_port, CEB => n105,
                           CK => clock, RB => resetn, Q => arx_r1_reg_13_port);
   arx_i1_reg_reg_6_inst : DFERPQ1 port map( D => data_in(6), CEB => n56, CK =>
                           clock, RB => resetn, Q => arx_i1_reg_6_port);
   arx_r3_reg_reg_12_inst : DFERPQ1 port map( D => a1_out_5_port, CEB => n1060,
                           CK => clock, RB => resetn, Q => arx_r3_reg_12_port);
   arx_r4_reg_reg_12_inst : DFERPQ1 port map( D => m3_out_12_port, CEB => n1070
                           , CK => clock, RB => resetn, Q => arx_r4_reg_12_port
                           );
   arx_r4_reg_reg_6_inst : DFERPQ1 port map( D => m3_out_6_port, CEB => n1070, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_6_port);
   arx_r2_reg_reg_12_inst : DFFRPQ1 port map( D => n80, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_12_port);
   arx_r1_reg_reg_12_inst : DFERPQ1 port map( D => m1_out_12_port, CEB => n105,
                           CK => clock, RB => resetn, Q => arx_r1_reg_12_port);
   arx_i1_reg_reg_5_inst : DFERPQ1 port map( D => data_in(5), CEB => n56, CK =>
                           clock, RB => resetn, Q => arx_i1_reg_5_port);
   arx_r3_reg_reg_11_inst : DFERPQ1 port map( D => a1_out_4_port, CEB => n1060,
                           CK => clock, RB => resetn, Q => arx_r3_reg_11_port);
   arx_r4_reg_reg_11_inst : DFERPQ1 port map( D => m3_out_11_port, CEB => n1070
                           , CK => clock, RB => resetn, Q => arx_r4_reg_11_port
                           );
   arx_r2_reg_reg_11_inst : DFFRPQ1 port map( D => n81, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_11_port);
   arx_r1_reg_reg_11_inst : DFERPQ1 port map( D => m1_out_11_port, CEB => n105,
                           CK => clock, RB => resetn, Q => arx_r1_reg_11_port);
   arx_i1_reg_reg_4_inst : DFERPQ1 port map( D => data_in(4), CEB => n56, CK =>
                           clock, RB => resetn, Q => arx_i1_reg_4_port);
   arx_r3_reg_reg_10_inst : DFERPQ1 port map( D => a1_out_3_port, CEB => n1060,
                           CK => clock, RB => resetn, Q => arx_r3_reg_10_port);
   arx_r4_reg_reg_10_inst : DFERPQ1 port map( D => m3_out_10_port, CEB => n1070
                           , CK => clock, RB => resetn, Q => arx_r4_reg_10_port
                           );
   arx_r2_reg_reg_10_inst : DFFRPQ1 port map( D => n82, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_10_port);
   arx_r1_reg_reg_10_inst : DFERPQ1 port map( D => m1_out_10_port, CEB => n105,
                           CK => clock, RB => resetn, Q => arx_r1_reg_10_port);
   arx_i1_reg_reg_3_inst : DFERPQ1 port map( D => data_in(3), CEB => n56, CK =>
                           clock, RB => resetn, Q => arx_i1_reg_3_port);
   arx_r3_reg_reg_9_inst : DFERPQ1 port map( D => a1_out_2_port, CEB => n1060, 
                           CK => clock, RB => resetn, Q => arx_r3_reg_9_port);
   arx_r4_reg_reg_9_inst : DFERPQ1 port map( D => m3_out_9_port, CEB => n1070, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_9_port);
   arx_r2_reg_reg_9_inst : DFFRPQ1 port map( D => n83, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_9_port);
   arx_r1_reg_reg_9_inst : DFERPQ1 port map( D => m1_out_9_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_9_port);
   arx_i1_reg_reg_2_inst : DFERPQ1 port map( D => data_in(2), CEB => n56, CK =>
                           clock, RB => resetn, Q => arx_i1_reg_2_port);
   arx_r3_reg_reg_8_inst : DFERPQ1 port map( D => a1_out_1_port, CEB => n1060, 
                           CK => clock, RB => resetn, Q => arx_r3_reg_8_port);
   arx_r4_reg_reg_8_inst : DFERPQ1 port map( D => m3_out_8_port, CEB => n1070, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_8_port);
   arx_r3_reg_reg_7_inst : DFERPQ1 port map( D => a1_out_0_port, CEB => n1060, 
                           CK => clock, RB => resetn, Q => arx_r3_reg_7_port);
   arx_r4_reg_reg_7_inst : DFERPQ1 port map( D => m3_out_7_port, CEB => n1070, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_7_port);
   arx_r2_reg_reg_8_inst : DFFRPQ1 port map( D => n84, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_8_port);
   arx_r1_reg_reg_8_inst : DFERPQ1 port map( D => m1_out_8_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_8_port);
   arx_i1_reg_reg_1_inst : DFERPQ1 port map( D => data_in(1), CEB => n56, CK =>
                           clock, RB => resetn, Q => arx_i1_reg_1_port);
   arx_r2_reg_reg_7_inst : DFFRPQ1 port map( D => n85, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_7_port);
   arx_r1_reg_reg_7_inst : DFERPQ1 port map( D => m1_out_7_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_7_port);
   arx_i1_reg_reg_0_inst : DFERPQ1 port map( D => data_in(0), CEB => n56, CK =>
                           clock, RB => resetn, Q => arx_i1_reg_0_port);
   arx_r1_reg_reg_6_inst : DFERPQ1 port map( D => m1_out_6_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_6_port);
   arx_r2_reg_reg_6_inst : DFFRPQ1 port map( D => n86, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_6_port);
   arx_r2_reg_reg_5_inst : DFFRPQ1 port map( D => n87, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_5_port);
   arx_r1_reg_reg_5_inst : DFERPQ1 port map( D => m1_out_5_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_5_port);
   arx_r2_reg_reg_4_inst : DFFRPQ1 port map( D => n88, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_4_port);
   arx_r1_reg_reg_4_inst : DFERPQ1 port map( D => m1_out_4_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_4_port);
   arx_d2_reg_reg_14_inst : DFERPQ1 port map( D => m1_in_r_7_port, CEB => n103,
                           CK => clock, RB => resetn, Q => m2_in_r_7_port);
   arx_d1_reg_reg_14_inst : DFERPQ1 port map( D => a1_out_7_port, CEB => n103, 
                           CK => clock, RB => resetn, Q => m1_in_r_7_port);
   arx_r2_reg_reg_3_inst : DFFRPQ1 port map( D => n89, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_3_port);
   arx_r1_reg_reg_3_inst : DFERPQ1 port map( D => m1_out_3_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_3_port);
   arx_d1_reg_reg_13_inst : DFERPQ1 port map( D => a1_out_6_port, CEB => n103, 
                           CK => clock, RB => resetn, Q => m1_in_r_6_port);
   arx_d1_reg_reg_12_inst : DFERPQ1 port map( D => a1_out_5_port, CEB => n102, 
                           CK => clock, RB => resetn, Q => m1_in_r_5_port);
   arx_d2_reg_reg_12_inst : DFERPQ1 port map( D => m1_in_r_5_port, CEB => n102,
                           CK => clock, RB => resetn, Q => m2_in_r_5_port);
   arx_d1_reg_reg_11_inst : DFERPQ1 port map( D => a1_out_4_port, CEB => n103, 
                           CK => clock, RB => resetn, Q => m1_in_r_4_port);
   arx_r2_reg_reg_2_inst : DFFRPQ1 port map( D => n90, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_2_port);
   arx_d2_reg_reg_13_inst : DFERPQ1 port map( D => m1_in_r_6_port, CEB => n55, 
                           CK => clock, RB => resetn, Q => m2_in_r_6_port);
   arx_r1_reg_reg_2_inst : DFERPQ1 port map( D => m1_out_2_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_2_port);
   arx_d1_reg_reg_10_inst : DFERPQ1 port map( D => a1_out_3_port, CEB => n102, 
                           CK => clock, RB => resetn, Q => m1_in_r_3_port);
   arx_d2_reg_reg_9_inst : DFERPQ1 port map( D => m1_in_r_2_port, CEB => n102, 
                           CK => clock, RB => resetn, Q => m2_in_r_2_port);
   arx_d2_reg_reg_11_inst : DFERPQ1 port map( D => m1_in_r_4_port, CEB => n103,
                           CK => clock, RB => resetn, Q => m2_in_r_4_port);
   arx_r1_reg_reg_0_inst : DFERPQ1 port map( D => m1_out_0_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_0_port);
   arx_r2_reg_reg_0_inst : DFFRPQ1 port map( D => n92, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_0_port);
   arx_d2_reg_reg_7_inst : DFERPQ1 port map( D => m1_in_r_0_port, CEB => n55, 
                           CK => clock, RB => resetn, Q => m2_in_r_0_port);
   arx_r1_reg_reg_1_inst : DFERPQ1 port map( D => m1_out_1_port, CEB => n105, 
                           CK => clock, RB => resetn, Q => arx_r1_reg_1_port);
   arx_d2_reg_reg_10_inst : DFERPQ1 port map( D => m1_in_r_3_port, CEB => n55, 
                           CK => clock, RB => resetn, Q => m2_in_r_3_port);
   arx_d1_reg_reg_9_inst : DFERPQ1 port map( D => a1_out_2_port, CEB => n103, 
                           CK => clock, RB => resetn, Q => m1_in_r_2_port);
   arx_d1_reg_reg_8_inst : DFERPQ1 port map( D => a1_out_1_port, CEB => n55, CK
                           => clock, RB => resetn, Q => m1_in_r_1_port);
   arx_d2_reg_reg_8_inst : DFERPQ1 port map( D => m1_in_r_1_port, CEB => n103, 
                           CK => clock, RB => resetn, Q => m2_in_r_1_port);
   arx_r2_reg_reg_1_inst : DFFRPQ1 port map( D => n91, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_1_port);
   arx_d1_reg_reg_7_inst : DFERPQ1 port map( D => a1_out_0_port, CEB => n102, 
                           CK => clock, RB => resetn, Q => m1_in_r_0_port);
   arx_state_reg_reg_1_inst : DFFRPQ1 port map( D => state_1_port, CK => clock,
                           RB => resetn, Q => arx_state_reg_1_port);
   arx_state_reg_reg_0_inst : DFFRPQ1 port map( D => n99, CK => clock, RB => 
                           resetn, Q => arx_state_reg_0_port);
   arx_o1_reg_reg_7_inst : DFERPQ1 port map( D => a2_out_7_port, CEB => n56, CK
                           => clock, RB => resetn, Q => data1_out(7));
   arx_o1_reg_reg_0_inst : DFERPQ1 port map( D => a2_out_0_port, CEB => n56, CK
                           => clock, RB => resetn, Q => data1_out(0));
   arx_o1_reg_reg_1_inst : DFERPQ1 port map( D => a2_out_1_port, CEB => n56, CK
                           => clock, RB => resetn, Q => data1_out(1));
   arx_o1_reg_reg_2_inst : DFERPQ1 port map( D => a2_out_2_port, CEB => n56, CK
                           => clock, RB => resetn, Q => data1_out(2));
   arx_o1_reg_reg_3_inst : DFERPQ1 port map( D => a2_out_3_port, CEB => n56, CK
                           => clock, RB => resetn, Q => data1_out(3));
   arx_o1_reg_reg_4_inst : DFERPQ1 port map( D => a2_out_4_port, CEB => n56, CK
                           => clock, RB => resetn, Q => data1_out(4));
   arx_o1_reg_reg_5_inst : DFERPQ1 port map( D => a2_out_5_port, CEB => n56, CK
                           => clock, RB => resetn, Q => data1_out(5));
   arx_o1_reg_reg_6_inst : DFERPQ1 port map( D => a2_out_6_port, CEB => n56, CK
                           => clock, RB => resetn, Q => data1_out(6));
   U135 : AND2D1 port map( A1 => arx_r1_reg_1_port, A2 => n99, Z => n93);
   U136 : AND2D1 port map( A1 => arx_r1_reg_0_port, A2 => n99, Z => n94);
   U137 : AND2D1 port map( A1 => arx_r1_reg_2_port, A2 => n99, Z => n95);
   U138 : AND2D1 port map( A1 => arx_r1_reg_3_port, A2 => n99, Z => n96);
   U139 : AND2D1 port map( A1 => arx_r1_reg_4_port, A2 => n99, Z => n97);
   U140 : AND2D1 port map( A1 => arx_r1_reg_6_port, A2 => n99, Z => n98);
   U141 : INVD1 port map( A => n57, Z => n1070);
   U142 : NOR2D1 port map( A1 => n1080, A2 => n99, Z => n57);
   U143 : OR2D1 port map( A1 => N137, A2 => n104, Z => n99);
   U144 : INVD1 port map( A => n100, Z => n104);
   U145 : INVD1 port map( A => N137, Z => n1060);
   U146 : NAN2D1 port map( A1 => n1060, A2 => n68, Z => m3_in_l_0);
   U147 : NAN2D1 port map( A1 => n102, A2 => n100, Z => m2_in_l_5_port);
   U148 : INVD1 port map( A => n55, Z => n1080);
   U149 : NOR2D1 port map( A1 => n57, A2 => n1170, Z => a1_in_r_14_port);
   U150 : NAN2M1D1 port map( A1 => state_1_port, A2 => n68, Z => n56);
   U151 : NAN2D1 port map( A1 => n103, A2 => n1060, Z => state_1_port);
   U152 : NAN2D1 port map( A1 => n55, A2 => n68, Z => n60);
   U153 : AND2D1 port map( A1 => arx_r2_reg_2_port, A2 => n1070, Z => 
                           a1_in_r_2_port);
   U154 : AND2D1 port map( A1 => arx_r2_reg_3_port, A2 => n1070, Z => 
                           a1_in_r_3_port);
   U155 : AND2D1 port map( A1 => arx_r2_reg_5_port, A2 => n1070, Z => 
                           a1_in_r_5_port);
   U156 : AND2D1 port map( A1 => arx_r2_reg_4_port, A2 => n1070, Z => 
                           a1_in_r_4_port);
   U157 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_7_port, B1 => n99, B2 
                           => arx_r1_reg_14_port, Z => a1_in_l_14_port);
   U158 : AND2D1 port map( A1 => arx_r2_reg_6_port, A2 => n1070, Z => 
                           a1_in_r_6_port);
   U159 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_0_port, B1 => n99, B2 
                           => arx_r1_reg_7_port, Z => a1_in_l_7_port);
   U160 : NOR2D1 port map( A1 => n57, A2 => n1100, Z => a1_in_r_7_port);
   U161 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_1_port, B1 => n99, B2 
                           => arx_r1_reg_8_port, Z => a1_in_l_8_port);
   U162 : NOR2D1 port map( A1 => n57, A2 => n1110, Z => a1_in_r_8_port);
   U163 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_2_port, B1 => n99, B2 
                           => arx_r1_reg_9_port, Z => a1_in_l_9_port);
   U164 : NOR2D1 port map( A1 => n57, A2 => n1120, Z => a1_in_r_9_port);
   U165 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_3_port, B1 => n99, B2 
                           => arx_r1_reg_10_port, Z => a1_in_l_10_port);
   U166 : NOR2D1 port map( A1 => n57, A2 => n1130, Z => a1_in_r_10_port);
   U167 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_4_port, B1 => n99, B2 
                           => arx_r1_reg_11_port, Z => a1_in_l_11_port);
   U168 : NOR2D1 port map( A1 => n57, A2 => n1140, Z => a1_in_r_11_port);
   U169 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_5_port, B1 => n99, B2 
                           => arx_r1_reg_12_port, Z => a1_in_l_12_port);
   U170 : NOR2D1 port map( A1 => n57, A2 => n1150, Z => a1_in_r_12_port);
   U171 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_6_port, B1 => n99, B2 
                           => arx_r1_reg_13_port, Z => a1_in_l_13_port);
   U172 : NOR2D1 port map( A1 => n57, A2 => n1160, Z => a1_in_r_13_port);
   U173 : AND2D1 port map( A1 => arx_r2_reg_1_port, A2 => n1070, Z => 
                           a1_in_r_1_port);
   U174 : OR2D1 port map( A1 => arx_state_reg_0_port, A2 => 
                           arx_state_reg_1_port, Z => n100);
   U175 : AND2D1 port map( A1 => arx_r2_reg_0_port, A2 => n1070, Z => 
                           a1_in_r_0_port);
   U176 : NOR2D1 port map( A1 => n1090, A2 => arx_state_reg_0_port, Z => N137);
   U177 : INVD1 port map( A => arx_state_reg_1_port, Z => n1090);
   U178 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => n1090, Z => n55);
   U179 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => 
                           arx_state_reg_1_port, Z => n68);
   U180 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => n1090, Z => n102);
   U181 : AND2D1 port map( A1 => m1_in_r_4_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_4_port);
   U182 : AND2D1 port map( A1 => m1_in_r_1_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_1_port);
   U183 : AND2D1 port map( A1 => m1_in_r_2_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_2_port);
   U184 : AND2D1 port map( A1 => m1_in_r_3_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_3_port);
   U185 : AND2D1 port map( A1 => m1_in_r_0_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_0_port);
   U186 : AND2D1 port map( A1 => m1_in_r_5_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_5_port);
   U187 : AND2D1 port map( A1 => arx_r1_reg_5_port, A2 => n99, Z => n101);
   U188 : AND2D1 port map( A1 => m1_in_r_6_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_6_port);
   U189 : AND2D1 port map( A1 => m1_in_r_7_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_7_port);
   U190 : AND2D1 port map( A1 => arx_r3_reg_9_port, A2 => n104, Z => 
                           a2_in_l_9_port);
   U191 : AND2D1 port map( A1 => arx_r4_reg_9_port, A2 => n104, Z => 
                           a2_in_r_9_port);
   U192 : AND2D1 port map( A1 => arx_r3_reg_10_port, A2 => n104, Z => 
                           a2_in_l_10_port);
   U193 : AND2D1 port map( A1 => arx_r4_reg_10_port, A2 => n104, Z => 
                           a2_in_r_10_port);
   U194 : AND2D1 port map( A1 => arx_r3_reg_11_port, A2 => n104, Z => 
                           a2_in_l_11_port);
   U195 : AND2D1 port map( A1 => arx_r4_reg_11_port, A2 => n104, Z => 
                           a2_in_r_11_port);
   U196 : AND2D1 port map( A1 => arx_r3_reg_12_port, A2 => n104, Z => 
                           a2_in_l_12_port);
   U197 : AND2D1 port map( A1 => arx_r4_reg_12_port, A2 => n104, Z => 
                           a2_in_r_12_port);
   U198 : AND2D1 port map( A1 => arx_r3_reg_13_port, A2 => n104, Z => 
                           a2_in_l_13_port);
   U199 : AND2D1 port map( A1 => arx_r4_reg_13_port, A2 => n104, Z => 
                           a2_in_r_13_port);
   U200 : AND2D1 port map( A1 => arx_r3_reg_8_port, A2 => n104, Z => 
                           a2_in_l_8_port);
   U201 : AND2D1 port map( A1 => arx_r4_reg_8_port, A2 => n104, Z => 
                           a2_in_r_8_port);
   U202 : AND2D1 port map( A1 => arx_r4_reg_7_port, A2 => n104, Z => 
                           a2_in_r_7_port);
   U203 : EXOR3D1 port map( A1 => a2_in_l_14_port, A2 => a2_in_r_14_port, A3 =>
                           add_224_carry_14_port, Z => N123);
   U204 : AND2D1 port map( A1 => arx_r3_reg_14_port, A2 => n104, Z => 
                           a2_in_l_14_port);
   U205 : AND2D1 port map( A1 => arx_r3_reg_7_port, A2 => n104, Z => 
                           a2_in_l_7_port);
   U206 : AO22D1 port map( A1 => arx_r2_reg_6_port, A2 => N137, B1 => 
                           m2_out_6_port, B2 => n60, Z => n86);
   U207 : AO22D1 port map( A1 => arx_r2_reg_5_port, A2 => N137, B1 => 
                           m2_out_5_port, B2 => n60, Z => n87);
   U208 : INVD1 port map( A => arx_r2_reg_7_port, Z => n1100);
   U209 : AO22D1 port map( A1 => arx_r2_reg_4_port, A2 => N137, B1 => 
                           m2_out_4_port, B2 => n60, Z => n88);
   U210 : INVD1 port map( A => arx_r2_reg_8_port, Z => n1110);
   U211 : AO22D1 port map( A1 => arx_r2_reg_3_port, A2 => N137, B1 => 
                           m2_out_3_port, B2 => n60, Z => n89);
   U212 : AND2D1 port map( A1 => arx_r4_reg_6_port, A2 => n104, Z => N115);
   U213 : INVD1 port map( A => arx_r2_reg_9_port, Z => n1120);
   U214 : AO22D1 port map( A1 => arx_r2_reg_2_port, A2 => N137, B1 => 
                           m2_out_2_port, B2 => n60, Z => n90);
   U215 : INVD1 port map( A => arx_r2_reg_10_port, Z => n1130);
   U216 : AO22D1 port map( A1 => arx_r2_reg_1_port, A2 => N137, B1 => 
                           m2_out_1_port, B2 => n60, Z => n91);
   U217 : INVD1 port map( A => arx_r2_reg_11_port, Z => n1140);
   U218 : AND2D1 port map( A1 => arx_r4_reg_14_port, A2 => n104, Z => 
                           a2_in_r_14_port);
   U219 : INVD1 port map( A => arx_r2_reg_12_port, Z => n1150);
   U220 : INVD1 port map( A => arx_r2_reg_13_port, Z => n1160);
   U221 : INVD1 port map( A => arx_r2_reg_14_port, Z => n1170);
   U222 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => n1090, Z => n103);
   U223 : AO22D1 port map( A1 => arx_r2_reg_0_port, A2 => N137, B1 => 
                           m2_out_0_port, B2 => n60, Z => n92);
   U224 : INVD1 port map( A => arx_state_reg_0_port, Z => n105);
   U225 : TIELO port map( Z => n1190);
   U226 : TIEHI port map( Z => n1180);
   U227 : EXOR2D1 port map( A1 => N123, A2 => add_416_C224_rn_carry_7_port, Z 
                           => a2_out_7_port);
   U228 : AND2D1 port map( A1 => add_416_C224_rn_carry_6_port, A2 => N122, Z =>
                           add_416_C224_rn_carry_7_port);
   U229 : EXOR2D1 port map( A1 => N122, A2 => add_416_C224_rn_carry_6_port, Z 
                           => a2_out_6_port);
   U230 : AND2D1 port map( A1 => add_416_C224_rn_carry_5_port, A2 => N121, Z =>
                           add_416_C224_rn_carry_6_port);
   U231 : EXOR2D1 port map( A1 => N121, A2 => add_416_C224_rn_carry_5_port, Z 
                           => a2_out_5_port);
   U232 : AND2D1 port map( A1 => add_416_C224_rn_carry_4_port, A2 => N120, Z =>
                           add_416_C224_rn_carry_5_port);
   U233 : EXOR2D1 port map( A1 => N120, A2 => add_416_C224_rn_carry_4_port, Z 
                           => a2_out_4_port);
   U234 : AND2D1 port map( A1 => add_416_C224_rn_carry_3_port, A2 => N119, Z =>
                           add_416_C224_rn_carry_4_port);
   U235 : EXOR2D1 port map( A1 => N119, A2 => add_416_C224_rn_carry_3_port, Z 
                           => a2_out_3_port);
   U236 : AND2D1 port map( A1 => add_416_C224_rn_carry_2_port, A2 => N118, Z =>
                           add_416_C224_rn_carry_3_port);
   U237 : EXOR2D1 port map( A1 => N118, A2 => add_416_C224_rn_carry_2_port, Z 
                           => a2_out_2_port);
   U238 : AND2D1 port map( A1 => add_416_C224_rn_carry_1_port, A2 => N117, Z =>
                           add_416_C224_rn_carry_2_port);
   U239 : EXOR2D1 port map( A1 => N117, A2 => add_416_C224_rn_carry_1_port, Z 
                           => a2_out_1_port);
   U240 : AND2D1 port map( A1 => N116, A2 => N115, Z => 
                           add_416_C224_rn_carry_1_port);
   U241 : EXOR2D1 port map( A1 => N115, A2 => N116, Z => a2_out_0_port);
   U242 : AND2D1 port map( A1 => a2_in_l_7_port, A2 => a2_in_r_7_port, Z => 
                           add_224_carry_8_port);
   U243 : EXOR2D1 port map( A1 => a2_in_r_7_port, A2 => a2_in_l_7_port, Z => 
                           N116);
   U244 : EXOR2D1 port map( A1 => N114, A2 => add_416_C223_rn_carry_7_port, Z 
                           => a1_out_7_port);
   U245 : AND2D1 port map( A1 => add_416_C223_rn_carry_6_port, A2 => N113, Z =>
                           add_416_C223_rn_carry_7_port);
   U246 : EXOR2D1 port map( A1 => N113, A2 => add_416_C223_rn_carry_6_port, Z 
                           => a1_out_6_port);
   U247 : AND2D1 port map( A1 => add_416_C223_rn_carry_5_port, A2 => N112, Z =>
                           add_416_C223_rn_carry_6_port);
   U248 : EXOR2D1 port map( A1 => N112, A2 => add_416_C223_rn_carry_5_port, Z 
                           => a1_out_5_port);
   U249 : AND2D1 port map( A1 => add_416_C223_rn_carry_4_port, A2 => N111, Z =>
                           add_416_C223_rn_carry_5_port);
   U250 : EXOR2D1 port map( A1 => N111, A2 => add_416_C223_rn_carry_4_port, Z 
                           => a1_out_4_port);
   U251 : AND2D1 port map( A1 => add_416_C223_rn_carry_3_port, A2 => N110, Z =>
                           add_416_C223_rn_carry_4_port);
   U252 : EXOR2D1 port map( A1 => N110, A2 => add_416_C223_rn_carry_3_port, Z 
                           => a1_out_3_port);
   U253 : AND2D1 port map( A1 => add_416_C223_rn_carry_2_port, A2 => N109, Z =>
                           add_416_C223_rn_carry_3_port);
   U254 : EXOR2D1 port map( A1 => N109, A2 => add_416_C223_rn_carry_2_port, Z 
                           => a1_out_2_port);
   U255 : AND2D1 port map( A1 => add_416_C223_rn_carry_1_port, A2 => N108, Z =>
                           add_416_C223_rn_carry_2_port);
   U256 : EXOR2D1 port map( A1 => N108, A2 => add_416_C223_rn_carry_1_port, Z 
                           => a1_out_1_port);
   U257 : AND2D1 port map( A1 => N107, A2 => N106, Z => 
                           add_416_C223_rn_carry_1_port);
   U258 : EXOR2D1 port map( A1 => N106, A2 => N107, Z => a1_out_0_port);

end hier_rtl_none_10;
