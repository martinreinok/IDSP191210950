
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_MAP1_overlapped is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type SIGNED is array (INTEGER range <>) of std_logic;

end CONV_PACK_MAP1_overlapped;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_MAP1_overlapped.all;

architecture flat_rtl_none_10 of MAP1_overlapped is

   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component MUXB2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIEHI
      port( Z : out std_logic);
   end component;
   
   component EXNOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2DL
      port( A0, A1, SL : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal arx_i1_reg_7_port, arx_i1_reg_6_port, arx_i1_reg_5_port, 
      arx_i1_reg_4_port, arx_i1_reg_3_port, arx_i1_reg_2_port, 
      arx_i1_reg_1_port, arx_i1_reg_0_port, arx_r1_reg_14_port, 
      arx_r1_reg_13_port, arx_r1_reg_12_port, arx_r1_reg_11_port, 
      arx_r1_reg_10_port, arx_r1_reg_9_port, arx_r1_reg_8_port, 
      arx_r1_reg_7_port, arx_r1_reg_6_port, arx_r1_reg_5_port, 
      arx_r1_reg_4_port, arx_r1_reg_3_port, arx_r1_reg_2_port, 
      arx_r1_reg_1_port, arx_r1_reg_0_port, arx_r2_reg_14_port, 
      arx_r2_reg_13_port, arx_r2_reg_12_port, arx_r2_reg_11_port, 
      arx_r2_reg_10_port, arx_r2_reg_9_port, arx_r2_reg_8_port, 
      arx_r2_reg_7_port, arx_r2_reg_6_port, arx_r2_reg_5_port, 
      arx_r2_reg_4_port, arx_r2_reg_3_port, arx_r2_reg_2_port, 
      arx_r2_reg_1_port, arx_r2_reg_0_port, arx_r3_reg_14_port, 
      arx_r3_reg_13_port, arx_r3_reg_12_port, arx_r3_reg_11_port, 
      arx_r3_reg_10_port, arx_r3_reg_9_port, arx_r3_reg_8_port, 
      arx_r3_reg_7_port, arx_r4_reg_14_port, arx_r4_reg_13_port, 
      arx_r4_reg_12_port, arx_r4_reg_11_port, arx_r4_reg_10_port, 
      arx_r4_reg_9_port, arx_r4_reg_8_port, arx_r4_reg_7_port, 
      arx_r4_reg_6_port, arx_state_reg_1_port, arx_state_reg_0_port, 
      m1_in_r_7_port, m1_in_r_6_port, m1_in_r_5_port, m1_in_r_4_port, 
      m1_in_r_3_port, m1_in_r_2_port, m1_in_r_1_port, m1_in_r_0_port, 
      m1_out_14_port, m1_out_13_port, m1_out_12_port, m1_out_11_port, 
      m1_out_10_port, m1_out_9_port, m1_out_8_port, m1_out_7_port, 
      m1_out_6_port, m1_out_5_port, m1_out_4_port, m1_out_3_port, m1_out_2_port
      , m1_out_1_port, m1_out_0_port, m2_in_l_5, m2_in_r_7_port, m2_in_r_6_port
      , m2_in_r_5_port, m2_in_r_4_port, m2_in_r_3_port, m2_in_r_2_port, 
      m2_in_r_1_port, m2_out_14_port, m2_out_13_port, m2_out_12_port, 
      m2_out_11_port, m2_out_10_port, m2_out_9_port, m2_out_8_port, 
      m2_out_7_port, m2_out_6_port, m2_out_5_port, m2_out_4_port, m2_out_3_port
      , m2_out_2_port, m2_out_1_port, m2_out_0_port, m3_in_l_0, m3_in_r_7_port,
      m3_in_r_6_port, m3_in_r_5_port, m3_in_r_4_port, m3_in_r_3_port, 
      m3_in_r_2_port, m3_in_r_1_port, m3_in_r_0_port, m3_out_15, m3_out_12_port
      , m3_out_11_port, m3_out_10_port, m3_out_9_port, m3_out_8_port, 
      m3_out_7_port, m3_out_6_port, a1_in_l_14_port, a1_in_l_13_port, 
      a1_in_l_12_port, a1_in_l_11_port, a1_in_l_10_port, a1_in_l_9_port, 
      a1_in_l_8_port, a1_in_l_7_port, a1_in_r_14_port, a1_in_r_13_port, 
      a1_in_r_12_port, a1_in_r_11_port, a1_in_r_10_port, a1_in_r_9_port, 
      a1_in_r_8_port, a1_in_r_7_port, a1_in_r_6_port, a1_in_r_5_port, 
      a1_in_r_4_port, a1_in_r_3_port, a1_in_r_2_port, a1_in_r_1_port, 
      a1_in_r_0_port, a1_out_7_port, a1_out_6_port, a1_out_5_port, 
      a1_out_4_port, a1_out_3_port, a1_out_2_port, a1_out_1_port, a1_out_0_port
      , a2_in_l_14_port, a2_in_l_13_port, a2_in_l_12_port, a2_in_l_11_port, 
      a2_in_l_10_port, a2_in_l_9_port, a2_in_l_8_port, a2_in_l_7_port, 
      a2_in_r_14_port, a2_in_r_13_port, a2_in_r_12_port, a2_in_r_11_port, 
      a2_in_r_10_port, a2_in_r_9_port, a2_in_r_8_port, a2_in_r_7_port, 
      a2_out_7_port, a2_out_6_port, a2_out_5_port, a2_out_4_port, a2_out_3_port
      , a2_out_2_port, a2_out_1_port, a2_out_0_port, state_1, N106, N107, N108,
      N109, N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, 
      N121, N122, N123, N137, n55, n56, n57, n58, n60, n61, n62, n63, n64, n65,
      n66, n67, n68, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89
      , n90, n91, n92, add_416_C224_rn_carry_1_port, 
      add_416_C224_rn_carry_2_port, add_416_C224_rn_carry_3_port, 
      add_416_C224_rn_carry_4_port, add_416_C224_rn_carry_5_port, 
      add_416_C224_rn_carry_6_port, add_416_C224_rn_carry_7_port, 
      add_224_carry_8_port, add_224_carry_9_port, add_224_carry_10_port, 
      add_224_carry_11_port, add_224_carry_12_port, add_224_carry_13_port, 
      add_224_carry_14_port, add_416_C223_rn_carry_1_port, 
      add_416_C223_rn_carry_2_port, add_416_C223_rn_carry_3_port, 
      add_416_C223_rn_carry_4_port, add_416_C223_rn_carry_5_port, 
      add_416_C223_rn_carry_6_port, add_416_C223_rn_carry_7_port, n93, n94, n95
      , n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n1060, n1070, 
      n1080, n1090, n1100, n1110, n1120, n1130, n1140, n1150, n1160, n1170, 
      n1180, n1190, n_1027, n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, 
      n_1034, n_1035, n_1036, n_1037, n_1038, n_1039, n_1040, n_1041, 
      add_223_n9, add_223_n8, add_223_n7, add_223_n6, add_223_n5, add_223_n4, 
      add_223_n3, add_223_n2, add_223_n1, add_223_carry_6_port, 
      add_223_carry_7_port, add_223_carry_8_port, add_223_carry_9_port, 
      add_223_carry_10_port, add_223_carry_11_port, add_223_carry_12_port, 
      add_223_carry_13_port, add_223_carry_14_port, mult_222_n_1011, 
      mult_222_n_1010, mult_222_n_1009, mult_222_n130, mult_222_n129, 
      mult_222_n128, mult_222_n127, mult_222_n126, mult_222_n125, mult_222_n124
      , mult_222_n123, mult_222_n122, mult_222_n121, mult_222_n119, 
      mult_222_n71, mult_222_n70, mult_222_n69, mult_222_n68, mult_222_n67, 
      mult_222_n66, mult_222_n65, mult_222_n64, mult_222_n63, mult_222_n62, 
      mult_222_n61, mult_222_n60, mult_222_n59, mult_222_n58, mult_222_n57, 
      mult_222_n56, mult_222_n55, mult_222_n54, mult_222_n53, mult_222_n52, 
      mult_222_n51, mult_222_n50, mult_222_n49, mult_222_n48, mult_222_n47, 
      mult_222_n46, mult_222_n45, mult_222_n44, mult_222_n43, mult_222_n42, 
      mult_222_n41, mult_222_n40, mult_222_n39, mult_222_n38, mult_222_n37, 
      mult_222_n36, mult_222_n35, mult_222_n33, mult_222_n32, mult_222_n31, 
      mult_222_n30, mult_222_n29, mult_222_n27, mult_222_n26, mult_222_n25, 
      mult_222_n24, mult_222_n23, mult_222_n21, mult_222_n20, mult_222_n19, 
      mult_222_n18, mult_222_n17, mult_222_n16, mult_222_n15, mult_222_n14, 
      mult_222_n13, mult_222_n12, mult_222_n11, mult_222_n10, mult_222_n9, 
      mult_222_n8, mult_222_n7, mult_222_n6, mult_222_n5, mult_222_n4, 
      mult_222_n3, mult_222_n2, mult_221_n212, mult_221_n211, mult_221_n210, 
      mult_221_n209, mult_221_n208, mult_221_n207, mult_221_n206, mult_221_n205
      , mult_221_n204, mult_221_n203, mult_221_n202, mult_221_n201, 
      mult_221_n200, mult_221_n199, mult_221_n198, mult_221_n197, mult_221_n196
      , mult_221_n195, mult_221_n194, mult_221_n193, mult_221_n192, 
      mult_221_n191, mult_221_n190, mult_221_n189, mult_221_n188, mult_221_n187
      , mult_221_n186, mult_221_n185, mult_221_n184, mult_221_n92, mult_221_n91
      , mult_221_n90, mult_221_n89, mult_221_n88, mult_221_n87, mult_221_n86, 
      mult_221_n83, mult_221_n82, mult_221_n81, mult_221_n80, mult_221_n79, 
      mult_221_n77, mult_221_n76, mult_221_n75, mult_221_n74, mult_221_n73, 
      mult_221_n72, mult_221_n71, mult_221_n70, mult_221_n69, mult_221_n68, 
      mult_221_n67, mult_221_n66, mult_221_n65, mult_221_n64, mult_221_n63, 
      mult_221_n62, mult_221_n60, mult_221_n57, mult_221_n56, mult_221_n55, 
      mult_221_n54, mult_221_n53, mult_221_n52, mult_221_n51, mult_221_n50, 
      mult_221_n48, mult_221_n47, mult_221_n46, mult_221_n45, mult_221_n44, 
      mult_221_n43, mult_221_n42, mult_221_n41, mult_221_n40, mult_221_n39, 
      mult_221_n38, mult_221_n37, mult_221_n36, mult_221_n35, mult_221_n34, 
      mult_221_n33, mult_221_n32, mult_221_n30, mult_221_n29, mult_221_n28, 
      mult_221_n27, mult_221_n26, mult_221_n25, mult_221_n24, mult_221_n23, 
      mult_221_n21, mult_221_n20, mult_221_n19, mult_221_n18, mult_221_n17, 
      mult_221_n16, mult_221_n14, mult_221_n12, mult_221_n11, mult_221_n10, 
      mult_221_n9, mult_221_n8, mult_221_n7, mult_221_n6, mult_221_n5, 
      mult_221_n4, mult_221_n3, mult_221_n2, mult_220_n187, mult_220_n186, 
      mult_220_n185, mult_220_n183, mult_220_n182, mult_220_n181, mult_220_n180
      , mult_220_n179, mult_220_n178, mult_220_n177, mult_220_n176, 
      mult_220_n175, mult_220_n174, mult_220_n126, mult_220_n112, mult_220_n111
      , mult_220_n110, mult_220_n109, mult_220_n108, mult_220_n107, 
      mult_220_n106, mult_220_n105, mult_220_n104, mult_220_n103, mult_220_n102
      , mult_220_n101, mult_220_n100, mult_220_n99, mult_220_n98, mult_220_n97,
      mult_220_n96, mult_220_n95, mult_220_n94, mult_220_n93, mult_220_n92, 
      mult_220_n91, mult_220_n90, mult_220_n89, mult_220_n88, mult_220_n87, 
      mult_220_n86, mult_220_n85, mult_220_n84, mult_220_n83, mult_220_n82, 
      mult_220_n62, mult_220_n61, mult_220_n60, mult_220_n59, mult_220_n58, 
      mult_220_n57, mult_220_n56, mult_220_n55, mult_220_n54, mult_220_n53, 
      mult_220_n52, mult_220_n51, mult_220_n50, mult_220_n49, mult_220_n48, 
      mult_220_n47, mult_220_n46, mult_220_n45, mult_220_n44, mult_220_n43, 
      mult_220_n42, mult_220_n41, mult_220_n40, mult_220_n39, mult_220_n37, 
      mult_220_n36, mult_220_n35, mult_220_n34, mult_220_n31, mult_220_n30, 
      mult_220_n29, mult_220_n28, mult_220_n27, mult_220_n26, mult_220_n25, 
      mult_220_n24, mult_220_n22, mult_220_n21, mult_220_n20, mult_220_n19, 
      mult_220_n18, mult_220_n16, mult_220_n15, mult_220_n14, mult_220_n13, 
      mult_220_n12, mult_220_n11, mult_220_n10, mult_220_n9, mult_220_n8, 
      mult_220_n7, mult_220_n6, mult_220_n5, mult_220_n4, mult_220_n3, 
      mult_220_n2 : std_logic;

begin
   
   U119 : OAI21D1 port map( A1 => n1060, A2 => n1170, B => n58, Z => n78);
   U120 : AOI22D1 port map( A1 => n104, A2 => a1_out_7_port, B1 => 
                           m2_out_14_port, B2 => n60, Z => n58);
   U121 : OAI21D1 port map( A1 => n1060, A2 => n1160, B => n61, Z => n79);
   U122 : AOI22D1 port map( A1 => n104, A2 => a1_out_6_port, B1 => 
                           m2_out_13_port, B2 => n60, Z => n61);
   U123 : OAI21D1 port map( A1 => n1060, A2 => n1150, B => n62, Z => n80);
   U124 : AOI22D1 port map( A1 => n104, A2 => a1_out_5_port, B1 => 
                           m2_out_12_port, B2 => n60, Z => n62);
   U125 : OAI21D1 port map( A1 => n1060, A2 => n1140, B => n63, Z => n81);
   U126 : AOI22D1 port map( A1 => n104, A2 => a1_out_4_port, B1 => 
                           m2_out_11_port, B2 => n60, Z => n63);
   U127 : OAI21D1 port map( A1 => n1060, A2 => n1130, B => n64, Z => n82);
   U128 : AOI22D1 port map( A1 => n104, A2 => a1_out_3_port, B1 => 
                           m2_out_10_port, B2 => n60, Z => n64);
   U129 : OAI21D1 port map( A1 => n1060, A2 => n1120, B => n65, Z => n83);
   U130 : AOI22D1 port map( A1 => n104, A2 => a1_out_2_port, B1 => 
                           m2_out_9_port, B2 => n60, Z => n65);
   U131 : OAI21D1 port map( A1 => n1060, A2 => n1110, B => n66, Z => n84);
   U132 : AOI22D1 port map( A1 => n104, A2 => a1_out_1_port, B1 => 
                           m2_out_8_port, B2 => n60, Z => n66);
   U133 : OAI21D1 port map( A1 => n1060, A2 => n1100, B => n67, Z => n85);
   U134 : AOI22D1 port map( A1 => n104, A2 => a1_out_0_port, B1 => 
                           m2_out_7_port, B2 => n60, Z => n67);
   add_224_U1_8 : ADFULD1 port map( A => a2_in_l_8_port, B => a2_in_r_8_port, 
                           CI => add_224_carry_8_port, CO => 
                           add_224_carry_9_port, S => N117);
   add_224_U1_9 : ADFULD1 port map( A => a2_in_l_9_port, B => a2_in_r_9_port, 
                           CI => add_224_carry_9_port, CO => 
                           add_224_carry_10_port, S => N118);
   add_224_U1_10 : ADFULD1 port map( A => a2_in_l_10_port, B => a2_in_r_10_port
                           , CI => add_224_carry_10_port, CO => 
                           add_224_carry_11_port, S => N119);
   add_224_U1_11 : ADFULD1 port map( A => a2_in_l_11_port, B => a2_in_r_11_port
                           , CI => add_224_carry_11_port, CO => 
                           add_224_carry_12_port, S => N120);
   add_224_U1_12 : ADFULD1 port map( A => a2_in_l_12_port, B => a2_in_r_12_port
                           , CI => add_224_carry_12_port, CO => 
                           add_224_carry_13_port, S => N121);
   add_224_U1_13 : ADFULD1 port map( A => a2_in_l_13_port, B => a2_in_r_13_port
                           , CI => add_224_carry_13_port, CO => 
                           add_224_carry_14_port, S => N122);
   arx_r3_reg_reg_14 : DFERPQ1 port map( D => a1_out_7_port, CEB => n1060, CK 
                           => clock, RB => resetn, Q => arx_r3_reg_14_port);
   arx_r4_reg_reg_14 : DFERPQ1 port map( D => m3_out_15, CEB => n1070, CK => 
                           clock, RB => resetn, Q => arx_r4_reg_14_port);
   arx_r2_reg_reg_14 : DFFRPQ1 port map( D => n78, CK => clock, RB => resetn, Q
                           => arx_r2_reg_14_port);
   arx_r1_reg_reg_14 : DFERPQ1 port map( D => m1_out_14_port, CEB => n105, CK 
                           => clock, RB => resetn, Q => arx_r1_reg_14_port);
   arx_i1_reg_reg_7 : DFERPQ1 port map( D => data_in(7), CEB => n56, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_7_port);
   arx_r3_reg_reg_13 : DFERPQ1 port map( D => a1_out_6_port, CEB => n1060, CK 
                           => clock, RB => resetn, Q => arx_r3_reg_13_port);
   arx_r4_reg_reg_13 : DFERPQ1 port map( D => m3_out_15, CEB => n1070, CK => 
                           clock, RB => resetn, Q => arx_r4_reg_13_port);
   arx_r2_reg_reg_13 : DFFRPQ1 port map( D => n79, CK => clock, RB => resetn, Q
                           => arx_r2_reg_13_port);
   arx_r1_reg_reg_13 : DFERPQ1 port map( D => m1_out_13_port, CEB => n105, CK 
                           => clock, RB => resetn, Q => arx_r1_reg_13_port);
   arx_i1_reg_reg_6 : DFERPQ1 port map( D => data_in(6), CEB => n56, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_6_port);
   arx_r3_reg_reg_12 : DFERPQ1 port map( D => a1_out_5_port, CEB => n1060, CK 
                           => clock, RB => resetn, Q => arx_r3_reg_12_port);
   arx_r4_reg_reg_12 : DFERPQ1 port map( D => m3_out_12_port, CEB => n1070, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_12_port);
   arx_r4_reg_reg_6 : DFERPQ1 port map( D => m3_out_6_port, CEB => n1070, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_6_port);
   arx_r2_reg_reg_12 : DFFRPQ1 port map( D => n80, CK => clock, RB => resetn, Q
                           => arx_r2_reg_12_port);
   arx_r1_reg_reg_12 : DFERPQ1 port map( D => m1_out_12_port, CEB => n105, CK 
                           => clock, RB => resetn, Q => arx_r1_reg_12_port);
   arx_i1_reg_reg_5 : DFERPQ1 port map( D => data_in(5), CEB => n56, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_5_port);
   arx_r3_reg_reg_11 : DFERPQ1 port map( D => a1_out_4_port, CEB => n1060, CK 
                           => clock, RB => resetn, Q => arx_r3_reg_11_port);
   arx_r4_reg_reg_11 : DFERPQ1 port map( D => m3_out_11_port, CEB => n1070, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_11_port);
   arx_r2_reg_reg_11 : DFFRPQ1 port map( D => n81, CK => clock, RB => resetn, Q
                           => arx_r2_reg_11_port);
   arx_r1_reg_reg_11 : DFERPQ1 port map( D => m1_out_11_port, CEB => n105, CK 
                           => clock, RB => resetn, Q => arx_r1_reg_11_port);
   arx_i1_reg_reg_4 : DFERPQ1 port map( D => data_in(4), CEB => n56, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_4_port);
   arx_r3_reg_reg_10 : DFERPQ1 port map( D => a1_out_3_port, CEB => n1060, CK 
                           => clock, RB => resetn, Q => arx_r3_reg_10_port);
   arx_r4_reg_reg_10 : DFERPQ1 port map( D => m3_out_10_port, CEB => n1070, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_10_port);
   arx_r2_reg_reg_10 : DFFRPQ1 port map( D => n82, CK => clock, RB => resetn, Q
                           => arx_r2_reg_10_port);
   arx_r1_reg_reg_10 : DFERPQ1 port map( D => m1_out_10_port, CEB => n105, CK 
                           => clock, RB => resetn, Q => arx_r1_reg_10_port);
   arx_i1_reg_reg_3 : DFERPQ1 port map( D => data_in(3), CEB => n56, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_3_port);
   arx_r3_reg_reg_9 : DFERPQ1 port map( D => a1_out_2_port, CEB => n1060, CK =>
                           clock, RB => resetn, Q => arx_r3_reg_9_port);
   arx_r4_reg_reg_9 : DFERPQ1 port map( D => m3_out_9_port, CEB => n1070, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_9_port);
   arx_r2_reg_reg_9 : DFFRPQ1 port map( D => n83, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_9_port);
   arx_r1_reg_reg_9 : DFERPQ1 port map( D => m1_out_9_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_9_port);
   arx_i1_reg_reg_2 : DFERPQ1 port map( D => data_in(2), CEB => n56, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_2_port);
   arx_r3_reg_reg_8 : DFERPQ1 port map( D => a1_out_1_port, CEB => n1060, CK =>
                           clock, RB => resetn, Q => arx_r3_reg_8_port);
   arx_r4_reg_reg_8 : DFERPQ1 port map( D => m3_out_8_port, CEB => n1070, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_8_port);
   arx_r3_reg_reg_7 : DFERPQ1 port map( D => a1_out_0_port, CEB => n1060, CK =>
                           clock, RB => resetn, Q => arx_r3_reg_7_port);
   arx_r4_reg_reg_7 : DFERPQ1 port map( D => m3_out_7_port, CEB => n1070, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_7_port);
   arx_r2_reg_reg_8 : DFFRPQ1 port map( D => n84, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_8_port);
   arx_r1_reg_reg_8 : DFERPQ1 port map( D => m1_out_8_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_8_port);
   arx_i1_reg_reg_1 : DFERPQ1 port map( D => data_in(1), CEB => n56, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_1_port);
   arx_r2_reg_reg_7 : DFFRPQ1 port map( D => n85, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_7_port);
   arx_r1_reg_reg_7 : DFERPQ1 port map( D => m1_out_7_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_7_port);
   arx_i1_reg_reg_0 : DFERPQ1 port map( D => data_in(0), CEB => n56, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_0_port);
   arx_r1_reg_reg_6 : DFERPQ1 port map( D => m1_out_6_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_6_port);
   arx_r2_reg_reg_6 : DFFRPQ1 port map( D => n86, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_6_port);
   arx_r2_reg_reg_5 : DFFRPQ1 port map( D => n87, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_5_port);
   arx_r1_reg_reg_5 : DFERPQ1 port map( D => m1_out_5_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_5_port);
   arx_r2_reg_reg_4 : DFFRPQ1 port map( D => n88, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_4_port);
   arx_r1_reg_reg_4 : DFERPQ1 port map( D => m1_out_4_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_4_port);
   arx_d2_reg_reg_14 : DFERPQ1 port map( D => m1_in_r_7_port, CEB => n103, CK 
                           => clock, RB => resetn, Q => m2_in_r_7_port);
   arx_d1_reg_reg_14 : DFERPQ1 port map( D => a1_out_7_port, CEB => n103, CK =>
                           clock, RB => resetn, Q => m1_in_r_7_port);
   arx_r2_reg_reg_3 : DFFRPQ1 port map( D => n89, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_3_port);
   arx_r1_reg_reg_3 : DFERPQ1 port map( D => m1_out_3_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_3_port);
   arx_d1_reg_reg_13 : DFERPQ1 port map( D => a1_out_6_port, CEB => n103, CK =>
                           clock, RB => resetn, Q => m1_in_r_6_port);
   arx_d1_reg_reg_12 : DFERPQ1 port map( D => a1_out_5_port, CEB => n102, CK =>
                           clock, RB => resetn, Q => m1_in_r_5_port);
   arx_d2_reg_reg_12 : DFERPQ1 port map( D => m1_in_r_5_port, CEB => n102, CK 
                           => clock, RB => resetn, Q => m2_in_r_5_port);
   arx_d1_reg_reg_11 : DFERPQ1 port map( D => a1_out_4_port, CEB => n103, CK =>
                           clock, RB => resetn, Q => m1_in_r_4_port);
   arx_r2_reg_reg_2 : DFFRPQ1 port map( D => n90, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_2_port);
   arx_d2_reg_reg_13 : DFERPQ1 port map( D => m1_in_r_6_port, CEB => n55, CK =>
                           clock, RB => resetn, Q => m2_in_r_6_port);
   arx_r1_reg_reg_2 : DFERPQ1 port map( D => m1_out_2_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_2_port);
   arx_d1_reg_reg_10 : DFERPQ1 port map( D => a1_out_3_port, CEB => n102, CK =>
                           clock, RB => resetn, Q => m1_in_r_3_port);
   arx_d2_reg_reg_9 : DFERPQ1 port map( D => m1_in_r_2_port, CEB => n102, CK =>
                           clock, RB => resetn, Q => m2_in_r_2_port);
   arx_d2_reg_reg_11 : DFERPQ1 port map( D => m1_in_r_4_port, CEB => n103, CK 
                           => clock, RB => resetn, Q => m2_in_r_4_port);
   arx_r1_reg_reg_0 : DFERPQ1 port map( D => m1_out_0_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_0_port);
   arx_r2_reg_reg_0 : DFFRPQ1 port map( D => n92, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_0_port);
   arx_d2_reg_reg_7 : DFERPQ1 port map( D => m1_in_r_0_port, CEB => n55, CK => 
                           clock, RB => resetn, Q => m2_out_0_port);
   arx_r1_reg_reg_1 : DFERPQ1 port map( D => m1_out_1_port, CEB => n105, CK => 
                           clock, RB => resetn, Q => arx_r1_reg_1_port);
   arx_d2_reg_reg_10 : DFERPQ1 port map( D => m1_in_r_3_port, CEB => n55, CK =>
                           clock, RB => resetn, Q => m2_in_r_3_port);
   arx_d1_reg_reg_9 : DFERPQ1 port map( D => a1_out_2_port, CEB => n103, CK => 
                           clock, RB => resetn, Q => m1_in_r_2_port);
   arx_d1_reg_reg_8 : DFERPQ1 port map( D => a1_out_1_port, CEB => n55, CK => 
                           clock, RB => resetn, Q => m1_in_r_1_port);
   arx_d2_reg_reg_8 : DFERPQ1 port map( D => m1_in_r_1_port, CEB => n103, CK =>
                           clock, RB => resetn, Q => m2_in_r_1_port);
   arx_r2_reg_reg_1 : DFFRPQ1 port map( D => n91, CK => clock, RB => resetn, Q 
                           => arx_r2_reg_1_port);
   arx_d1_reg_reg_7 : DFERPQ1 port map( D => a1_out_0_port, CEB => n102, CK => 
                           clock, RB => resetn, Q => m1_in_r_0_port);
   arx_state_reg_reg_1 : DFFRPQ1 port map( D => state_1, CK => clock, RB => 
                           resetn, Q => arx_state_reg_1_port);
   arx_state_reg_reg_0 : DFFRPQ1 port map( D => n99, CK => clock, RB => resetn,
                           Q => arx_state_reg_0_port);
   arx_o1_reg_reg_7 : DFERPQ1 port map( D => a2_out_7_port, CEB => n56, CK => 
                           clock, RB => resetn, Q => data1_out(7));
   arx_o1_reg_reg_0 : DFERPQ1 port map( D => a2_out_0_port, CEB => n56, CK => 
                           clock, RB => resetn, Q => data1_out(0));
   arx_o1_reg_reg_1 : DFERPQ1 port map( D => a2_out_1_port, CEB => n56, CK => 
                           clock, RB => resetn, Q => data1_out(1));
   arx_o1_reg_reg_2 : DFERPQ1 port map( D => a2_out_2_port, CEB => n56, CK => 
                           clock, RB => resetn, Q => data1_out(2));
   arx_o1_reg_reg_3 : DFERPQ1 port map( D => a2_out_3_port, CEB => n56, CK => 
                           clock, RB => resetn, Q => data1_out(3));
   arx_o1_reg_reg_4 : DFERPQ1 port map( D => a2_out_4_port, CEB => n56, CK => 
                           clock, RB => resetn, Q => data1_out(4));
   arx_o1_reg_reg_5 : DFERPQ1 port map( D => a2_out_5_port, CEB => n56, CK => 
                           clock, RB => resetn, Q => data1_out(5));
   arx_o1_reg_reg_6 : DFERPQ1 port map( D => a2_out_6_port, CEB => n56, CK => 
                           clock, RB => resetn, Q => data1_out(6));
   U135 : AND2D1 port map( A1 => arx_r1_reg_1_port, A2 => n99, Z => n93);
   U136 : AND2D1 port map( A1 => arx_r1_reg_0_port, A2 => n99, Z => n94);
   U137 : AND2D1 port map( A1 => arx_r1_reg_2_port, A2 => n99, Z => n95);
   U138 : AND2D1 port map( A1 => arx_r1_reg_3_port, A2 => n99, Z => n96);
   U139 : AND2D1 port map( A1 => arx_r1_reg_4_port, A2 => n99, Z => n97);
   U140 : AND2D1 port map( A1 => arx_r1_reg_6_port, A2 => n99, Z => n98);
   U141 : INVD1 port map( A => n57, Z => n1070);
   U142 : NOR2D1 port map( A1 => n1080, A2 => n99, Z => n57);
   U143 : OR2D1 port map( A1 => N137, A2 => n104, Z => n99);
   U144 : INVD1 port map( A => n100, Z => n104);
   U145 : INVD1 port map( A => N137, Z => n1060);
   U146 : NAN2D1 port map( A1 => n1060, A2 => n68, Z => m3_in_l_0);
   U147 : NAN2D1 port map( A1 => n102, A2 => n100, Z => m2_in_l_5);
   U148 : INVD1 port map( A => n55, Z => n1080);
   U149 : NOR2D1 port map( A1 => n57, A2 => n1170, Z => a1_in_r_14_port);
   U150 : NAN2M1D1 port map( A1 => state_1, A2 => n68, Z => n56);
   U151 : NAN2D1 port map( A1 => n103, A2 => n1060, Z => state_1);
   U152 : NAN2D1 port map( A1 => n55, A2 => n68, Z => n60);
   U153 : AND2D1 port map( A1 => arx_r2_reg_2_port, A2 => n1070, Z => 
                           a1_in_r_2_port);
   U154 : AND2D1 port map( A1 => arx_r2_reg_3_port, A2 => n1070, Z => 
                           a1_in_r_3_port);
   U155 : AND2D1 port map( A1 => arx_r2_reg_5_port, A2 => n1070, Z => 
                           a1_in_r_5_port);
   U156 : AND2D1 port map( A1 => arx_r2_reg_4_port, A2 => n1070, Z => 
                           a1_in_r_4_port);
   U157 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_7_port, B1 => n99, B2 
                           => arx_r1_reg_14_port, Z => a1_in_l_14_port);
   U158 : AND2D1 port map( A1 => arx_r2_reg_6_port, A2 => n1070, Z => 
                           a1_in_r_6_port);
   U159 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_0_port, B1 => n99, B2 
                           => arx_r1_reg_7_port, Z => a1_in_l_7_port);
   U160 : NOR2D1 port map( A1 => n57, A2 => n1100, Z => a1_in_r_7_port);
   U161 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_1_port, B1 => n99, B2 
                           => arx_r1_reg_8_port, Z => a1_in_l_8_port);
   U162 : NOR2D1 port map( A1 => n57, A2 => n1110, Z => a1_in_r_8_port);
   U163 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_2_port, B1 => n99, B2 
                           => arx_r1_reg_9_port, Z => a1_in_l_9_port);
   U164 : NOR2D1 port map( A1 => n57, A2 => n1120, Z => a1_in_r_9_port);
   U165 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_3_port, B1 => n99, B2 
                           => arx_r1_reg_10_port, Z => a1_in_l_10_port);
   U166 : NOR2D1 port map( A1 => n57, A2 => n1130, Z => a1_in_r_10_port);
   U167 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_4_port, B1 => n99, B2 
                           => arx_r1_reg_11_port, Z => a1_in_l_11_port);
   U168 : NOR2D1 port map( A1 => n57, A2 => n1140, Z => a1_in_r_11_port);
   U169 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_5_port, B1 => n99, B2 
                           => arx_r1_reg_12_port, Z => a1_in_l_12_port);
   U170 : NOR2D1 port map( A1 => n57, A2 => n1150, Z => a1_in_r_12_port);
   U171 : AO22D1 port map( A1 => n1080, A2 => arx_i1_reg_6_port, B1 => n99, B2 
                           => arx_r1_reg_13_port, Z => a1_in_l_13_port);
   U172 : NOR2D1 port map( A1 => n57, A2 => n1160, Z => a1_in_r_13_port);
   U173 : AND2D1 port map( A1 => arx_r2_reg_1_port, A2 => n1070, Z => 
                           a1_in_r_1_port);
   U174 : OR2D1 port map( A1 => arx_state_reg_0_port, A2 => 
                           arx_state_reg_1_port, Z => n100);
   U175 : AND2D1 port map( A1 => arx_r2_reg_0_port, A2 => n1070, Z => 
                           a1_in_r_0_port);
   U176 : NOR2D1 port map( A1 => n1090, A2 => arx_state_reg_0_port, Z => N137);
   U177 : INVD1 port map( A => arx_state_reg_1_port, Z => n1090);
   U178 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => n1090, Z => n55);
   U179 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => 
                           arx_state_reg_1_port, Z => n68);
   U180 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => n1090, Z => n102);
   U181 : AND2D1 port map( A1 => m1_in_r_4_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_4_port);
   U182 : AND2D1 port map( A1 => m1_in_r_1_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_1_port);
   U183 : AND2D1 port map( A1 => m1_in_r_2_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_2_port);
   U184 : AND2D1 port map( A1 => m1_in_r_3_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_3_port);
   U185 : AND2D1 port map( A1 => m1_in_r_0_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_0_port);
   U186 : AND2D1 port map( A1 => m1_in_r_5_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_5_port);
   U187 : AND2D1 port map( A1 => arx_r1_reg_5_port, A2 => n99, Z => n101);
   U188 : AND2D1 port map( A1 => m1_in_r_6_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_6_port);
   U189 : AND2D1 port map( A1 => m1_in_r_7_port, A2 => m3_in_l_0, Z => 
                           m3_in_r_7_port);
   U190 : AND2D1 port map( A1 => arx_r3_reg_9_port, A2 => n104, Z => 
                           a2_in_l_9_port);
   U191 : AND2D1 port map( A1 => arx_r4_reg_9_port, A2 => n104, Z => 
                           a2_in_r_9_port);
   U192 : AND2D1 port map( A1 => arx_r3_reg_10_port, A2 => n104, Z => 
                           a2_in_l_10_port);
   U193 : AND2D1 port map( A1 => arx_r4_reg_10_port, A2 => n104, Z => 
                           a2_in_r_10_port);
   U194 : AND2D1 port map( A1 => arx_r3_reg_11_port, A2 => n104, Z => 
                           a2_in_l_11_port);
   U195 : AND2D1 port map( A1 => arx_r4_reg_11_port, A2 => n104, Z => 
                           a2_in_r_11_port);
   U196 : AND2D1 port map( A1 => arx_r3_reg_12_port, A2 => n104, Z => 
                           a2_in_l_12_port);
   U197 : AND2D1 port map( A1 => arx_r4_reg_12_port, A2 => n104, Z => 
                           a2_in_r_12_port);
   U198 : AND2D1 port map( A1 => arx_r3_reg_13_port, A2 => n104, Z => 
                           a2_in_l_13_port);
   U199 : AND2D1 port map( A1 => arx_r4_reg_13_port, A2 => n104, Z => 
                           a2_in_r_13_port);
   U200 : AND2D1 port map( A1 => arx_r3_reg_8_port, A2 => n104, Z => 
                           a2_in_l_8_port);
   U201 : AND2D1 port map( A1 => arx_r4_reg_8_port, A2 => n104, Z => 
                           a2_in_r_8_port);
   U202 : AND2D1 port map( A1 => arx_r4_reg_7_port, A2 => n104, Z => 
                           a2_in_r_7_port);
   U203 : EXOR3D1 port map( A1 => a2_in_l_14_port, A2 => a2_in_r_14_port, A3 =>
                           add_224_carry_14_port, Z => N123);
   U204 : AND2D1 port map( A1 => arx_r3_reg_14_port, A2 => n104, Z => 
                           a2_in_l_14_port);
   U205 : AND2D1 port map( A1 => arx_r3_reg_7_port, A2 => n104, Z => 
                           a2_in_l_7_port);
   U206 : AO22D1 port map( A1 => arx_r2_reg_6_port, A2 => N137, B1 => 
                           m2_out_6_port, B2 => n60, Z => n86);
   U207 : AO22D1 port map( A1 => arx_r2_reg_5_port, A2 => N137, B1 => 
                           m2_out_5_port, B2 => n60, Z => n87);
   U208 : INVD1 port map( A => arx_r2_reg_7_port, Z => n1100);
   U209 : AO22D1 port map( A1 => arx_r2_reg_4_port, A2 => N137, B1 => 
                           m2_out_4_port, B2 => n60, Z => n88);
   U210 : INVD1 port map( A => arx_r2_reg_8_port, Z => n1110);
   U211 : AO22D1 port map( A1 => arx_r2_reg_3_port, A2 => N137, B1 => 
                           m2_out_3_port, B2 => n60, Z => n89);
   U212 : AND2D1 port map( A1 => arx_r4_reg_6_port, A2 => n104, Z => N115);
   U213 : INVD1 port map( A => arx_r2_reg_9_port, Z => n1120);
   U214 : AO22D1 port map( A1 => arx_r2_reg_2_port, A2 => N137, B1 => 
                           m2_out_2_port, B2 => n60, Z => n90);
   U215 : INVD1 port map( A => arx_r2_reg_10_port, Z => n1130);
   U216 : AO22D1 port map( A1 => arx_r2_reg_1_port, A2 => N137, B1 => 
                           m2_out_1_port, B2 => n60, Z => n91);
   U217 : INVD1 port map( A => arx_r2_reg_11_port, Z => n1140);
   U218 : AND2D1 port map( A1 => arx_r4_reg_14_port, A2 => n104, Z => 
                           a2_in_r_14_port);
   U219 : INVD1 port map( A => arx_r2_reg_12_port, Z => n1150);
   U220 : INVD1 port map( A => arx_r2_reg_13_port, Z => n1160);
   U221 : INVD1 port map( A => arx_r2_reg_14_port, Z => n1170);
   U222 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => n1090, Z => n103);
   U223 : AO22D1 port map( A1 => arx_r2_reg_0_port, A2 => N137, B1 => 
                           m2_out_0_port, B2 => n60, Z => n92);
   U224 : INVD1 port map( A => arx_state_reg_0_port, Z => n105);
   U225 : TIELO port map( Z => n1190);
   U226 : TIEHI port map( Z => n1180);
   U227 : EXOR2D1 port map( A1 => N123, A2 => add_416_C224_rn_carry_7_port, Z 
                           => a2_out_7_port);
   U228 : AND2D1 port map( A1 => add_416_C224_rn_carry_6_port, A2 => N122, Z =>
                           add_416_C224_rn_carry_7_port);
   U229 : EXOR2D1 port map( A1 => N122, A2 => add_416_C224_rn_carry_6_port, Z 
                           => a2_out_6_port);
   U230 : AND2D1 port map( A1 => add_416_C224_rn_carry_5_port, A2 => N121, Z =>
                           add_416_C224_rn_carry_6_port);
   U231 : EXOR2D1 port map( A1 => N121, A2 => add_416_C224_rn_carry_5_port, Z 
                           => a2_out_5_port);
   U232 : AND2D1 port map( A1 => add_416_C224_rn_carry_4_port, A2 => N120, Z =>
                           add_416_C224_rn_carry_5_port);
   U233 : EXOR2D1 port map( A1 => N120, A2 => add_416_C224_rn_carry_4_port, Z 
                           => a2_out_4_port);
   U234 : AND2D1 port map( A1 => add_416_C224_rn_carry_3_port, A2 => N119, Z =>
                           add_416_C224_rn_carry_4_port);
   U235 : EXOR2D1 port map( A1 => N119, A2 => add_416_C224_rn_carry_3_port, Z 
                           => a2_out_3_port);
   U236 : AND2D1 port map( A1 => add_416_C224_rn_carry_2_port, A2 => N118, Z =>
                           add_416_C224_rn_carry_3_port);
   U237 : EXOR2D1 port map( A1 => N118, A2 => add_416_C224_rn_carry_2_port, Z 
                           => a2_out_2_port);
   U238 : AND2D1 port map( A1 => add_416_C224_rn_carry_1_port, A2 => N117, Z =>
                           add_416_C224_rn_carry_2_port);
   U239 : EXOR2D1 port map( A1 => N117, A2 => add_416_C224_rn_carry_1_port, Z 
                           => a2_out_1_port);
   U240 : AND2D1 port map( A1 => N116, A2 => N115, Z => 
                           add_416_C224_rn_carry_1_port);
   U241 : EXOR2D1 port map( A1 => N115, A2 => N116, Z => a2_out_0_port);
   U242 : AND2D1 port map( A1 => a2_in_l_7_port, A2 => a2_in_r_7_port, Z => 
                           add_224_carry_8_port);
   U243 : EXOR2D1 port map( A1 => a2_in_r_7_port, A2 => a2_in_l_7_port, Z => 
                           N116);
   U244 : EXOR2D1 port map( A1 => N114, A2 => add_416_C223_rn_carry_7_port, Z 
                           => a1_out_7_port);
   U245 : AND2D1 port map( A1 => add_416_C223_rn_carry_6_port, A2 => N113, Z =>
                           add_416_C223_rn_carry_7_port);
   U246 : EXOR2D1 port map( A1 => N113, A2 => add_416_C223_rn_carry_6_port, Z 
                           => a1_out_6_port);
   U247 : AND2D1 port map( A1 => add_416_C223_rn_carry_5_port, A2 => N112, Z =>
                           add_416_C223_rn_carry_6_port);
   U248 : EXOR2D1 port map( A1 => N112, A2 => add_416_C223_rn_carry_5_port, Z 
                           => a1_out_5_port);
   U249 : AND2D1 port map( A1 => add_416_C223_rn_carry_4_port, A2 => N111, Z =>
                           add_416_C223_rn_carry_5_port);
   U250 : EXOR2D1 port map( A1 => N111, A2 => add_416_C223_rn_carry_4_port, Z 
                           => a1_out_4_port);
   U251 : AND2D1 port map( A1 => add_416_C223_rn_carry_3_port, A2 => N110, Z =>
                           add_416_C223_rn_carry_4_port);
   U252 : EXOR2D1 port map( A1 => N110, A2 => add_416_C223_rn_carry_3_port, Z 
                           => a1_out_3_port);
   U253 : AND2D1 port map( A1 => add_416_C223_rn_carry_2_port, A2 => N109, Z =>
                           add_416_C223_rn_carry_3_port);
   U254 : EXOR2D1 port map( A1 => N109, A2 => add_416_C223_rn_carry_2_port, Z 
                           => a1_out_2_port);
   U255 : AND2D1 port map( A1 => add_416_C223_rn_carry_1_port, A2 => N108, Z =>
                           add_416_C223_rn_carry_2_port);
   U256 : EXOR2D1 port map( A1 => N108, A2 => add_416_C223_rn_carry_1_port, Z 
                           => a1_out_1_port);
   U257 : AND2D1 port map( A1 => N107, A2 => N106, Z => 
                           add_416_C223_rn_carry_1_port);
   U258 : EXOR2D1 port map( A1 => N106, A2 => N107, Z => a1_out_0_port);
   add_223_U10 : OAI211D1 port map( A1 => n93, A2 => a1_in_r_1_port, B => n94, 
                           C => a1_in_r_0_port, Z => add_223_n9);
   add_223_U9 : OAI21M20D1 port map( A1 => n93, A2 => a1_in_r_1_port, B => 
                           add_223_n9, Z => add_223_n7);
   add_223_U8 : OAI21D1 port map( A1 => n95, A2 => add_223_n7, B => 
                           a1_in_r_2_port, Z => add_223_n8);
   add_223_U7 : OAI21M20D1 port map( A1 => add_223_n7, A2 => n95, B => 
                           add_223_n8, Z => add_223_n5);
   add_223_U6 : OAI21D1 port map( A1 => n96, A2 => add_223_n5, B => 
                           a1_in_r_3_port, Z => add_223_n6);
   add_223_U5 : OAI21M20D1 port map( A1 => add_223_n5, A2 => n96, B => 
                           add_223_n6, Z => add_223_n3);
   add_223_U4 : OAI21D1 port map( A1 => n97, A2 => add_223_n3, B => 
                           a1_in_r_4_port, Z => add_223_n4);
   add_223_U3 : OAI21M20D1 port map( A1 => add_223_n3, A2 => n97, B => 
                           add_223_n4, Z => add_223_n1);
   add_223_U2 : OAI21D1 port map( A1 => n101, A2 => add_223_n1, B => 
                           a1_in_r_5_port, Z => add_223_n2);
   add_223_U1 : OAI21M20D1 port map( A1 => add_223_n1, A2 => n101, B => 
                           add_223_n2, Z => add_223_carry_6_port);
   add_223_U1_14 : EXOR3D1 port map( A1 => a1_in_l_14_port, A2 => 
                           a1_in_r_14_port, A3 => add_223_carry_14_port, Z => 
                           N114);
   add_223_U1_6 : ADFULD1 port map( A => n98, B => a1_in_r_6_port, CI => 
                           add_223_carry_6_port, CO => add_223_carry_7_port, S 
                           => N106);
   add_223_U1_7 : ADFULD1 port map( A => a1_in_l_7_port, B => a1_in_r_7_port, 
                           CI => add_223_carry_7_port, CO => 
                           add_223_carry_8_port, S => N107);
   add_223_U1_8 : ADFULD1 port map( A => a1_in_l_8_port, B => a1_in_r_8_port, 
                           CI => add_223_carry_8_port, CO => 
                           add_223_carry_9_port, S => N108);
   add_223_U1_9 : ADFULD1 port map( A => a1_in_l_9_port, B => a1_in_r_9_port, 
                           CI => add_223_carry_9_port, CO => 
                           add_223_carry_10_port, S => N109);
   add_223_U1_10 : ADFULD1 port map( A => a1_in_l_10_port, B => a1_in_r_10_port
                           , CI => add_223_carry_10_port, CO => 
                           add_223_carry_11_port, S => N110);
   add_223_U1_11 : ADFULD1 port map( A => a1_in_l_11_port, B => a1_in_r_11_port
                           , CI => add_223_carry_11_port, CO => 
                           add_223_carry_12_port, S => N111);
   add_223_U1_12 : ADFULD1 port map( A => a1_in_l_12_port, B => a1_in_r_12_port
                           , CI => add_223_carry_12_port, CO => 
                           add_223_carry_13_port, S => N112);
   add_223_U1_13 : ADFULD1 port map( A => a1_in_l_13_port, B => a1_in_r_13_port
                           , CI => add_223_carry_13_port, CO => 
                           add_223_carry_14_port, S => N113);
   mult_222_U118 : NAN2D1 port map( A1 => m3_in_l_0, A2 => m3_in_r_4_port, Z =>
                           mult_222_n23);
   mult_222_U117 : NAN2D1 port map( A1 => m3_in_l_0, A2 => m3_in_r_3_port, Z =>
                           mult_222_n29);
   mult_222_U116 : NAN2D1 port map( A1 => m3_in_l_0, A2 => m3_in_r_2_port, Z =>
                           mult_222_n35);
   mult_222_U115 : NAN2D1 port map( A1 => m3_in_l_0, A2 => m3_in_r_7_port, Z =>
                           mult_222_n46);
   mult_222_U114 : NOR2D1 port map( A1 => mult_222_n121, A2 => mult_222_n119, Z
                           => mult_222_n47);
   mult_222_U113 : NOR2D1 port map( A1 => mult_222_n122, A2 => mult_222_n119, Z
                           => mult_222_n48);
   mult_222_U112 : NOR2D1 port map( A1 => mult_222_n129, A2 => mult_222_n119, Z
                           => mult_222_n49);
   mult_222_U111 : NOR2D1 port map( A1 => mult_222_n130, A2 => mult_222_n119, Z
                           => mult_222_n50);
   mult_222_U110 : NAN2D1 port map( A1 => m3_in_l_0, A2 => m3_in_r_7_port, Z =>
                           mult_222_n51);
   mult_222_U109 : NOR2D1 port map( A1 => mult_222_n121, A2 => mult_222_n119, Z
                           => mult_222_n52);
   mult_222_U108 : NOR2D1 port map( A1 => mult_222_n122, A2 => mult_222_n119, Z
                           => mult_222_n53);
   mult_222_U107 : NOR2D1 port map( A1 => mult_222_n123, A2 => mult_222_n119, Z
                           => mult_222_n54);
   mult_222_U106 : NOR2D1 port map( A1 => mult_222_n125, A2 => mult_222_n119, Z
                           => mult_222_n55);
   mult_222_U105 : NOR2D1 port map( A1 => mult_222_n127, A2 => mult_222_n119, Z
                           => mult_222_n56);
   mult_222_U104 : NOR2D1 port map( A1 => mult_222_n129, A2 => mult_222_n119, Z
                           => mult_222_n57);
   mult_222_U103 : NOR2D1 port map( A1 => mult_222_n130, A2 => mult_222_n119, Z
                           => mult_222_n58);
   mult_222_U102 : NAN2D1 port map( A1 => m3_in_l_0, A2 => m3_in_r_7_port, Z =>
                           mult_222_n59);
   mult_222_U101 : NOR2D1 port map( A1 => mult_222_n121, A2 => mult_222_n119, Z
                           => mult_222_n60);
   mult_222_U100 : NOR2D1 port map( A1 => mult_222_n122, A2 => mult_222_n119, Z
                           => mult_222_n61);
   mult_222_U99 : NOR2D1 port map( A1 => mult_222_n123, A2 => mult_222_n119, Z 
                           => mult_222_n62);
   mult_222_U98 : NOR2D1 port map( A1 => mult_222_n125, A2 => mult_222_n119, Z 
                           => mult_222_n63);
   mult_222_U97 : NOR2D1 port map( A1 => mult_222_n127, A2 => mult_222_n119, Z 
                           => mult_222_n64);
   mult_222_U96 : NOR2D1 port map( A1 => mult_222_n129, A2 => mult_222_n119, Z 
                           => mult_222_n65);
   mult_222_U95 : NOR2D1 port map( A1 => mult_222_n130, A2 => mult_222_n119, Z 
                           => mult_222_n66);
   mult_222_U94 : NAN2D1 port map( A1 => m3_in_r_7_port, A2 => m3_in_l_0, Z => 
                           mult_222_n67);
   mult_222_U93 : NOR2D1 port map( A1 => mult_222_n119, A2 => mult_222_n121, Z 
                           => mult_222_n68);
   mult_222_U92 : NOR2D1 port map( A1 => mult_222_n119, A2 => mult_222_n122, Z 
                           => mult_222_n69);
   mult_222_U91 : NOR2D1 port map( A1 => mult_222_n119, A2 => mult_222_n123, Z 
                           => mult_222_n70);
   mult_222_U90 : NOR2D1 port map( A1 => mult_222_n119, A2 => mult_222_n125, Z 
                           => mult_222_n71);
   mult_222_U89 : INVD1 port map( A => m3_in_r_6_port, Z => mult_222_n121);
   mult_222_U88 : INVD1 port map( A => m3_in_r_5_port, Z => mult_222_n122);
   mult_222_U87 : INVD1 port map( A => m3_in_r_0_port, Z => mult_222_n130);
   mult_222_U86 : INVD1 port map( A => m3_in_r_1_port, Z => mult_222_n129);
   mult_222_U85 : INVD1 port map( A => mult_222_n23, Z => mult_222_n124);
   mult_222_U84 : INVD1 port map( A => mult_222_n29, Z => mult_222_n126);
   mult_222_U83 : INVD1 port map( A => mult_222_n35, Z => mult_222_n128);
   mult_222_U82 : INVD1 port map( A => m3_in_r_3_port, Z => mult_222_n125);
   mult_222_U81 : INVD1 port map( A => m3_in_r_2_port, Z => mult_222_n127);
   mult_222_U80 : INVD1 port map( A => m3_in_r_4_port, Z => mult_222_n123);
   mult_222_U79 : INVD1 port map( A => mult_222_n2, Z => m3_out_15);
   mult_222_U78 : INVD1 port map( A => m3_in_l_0, Z => mult_222_n119);
   mult_222_U30 : ADHALFDL port map( A => mult_222_n65, B => mult_222_n70, CO 
                           => mult_222_n44, S => mult_222_n45);
   mult_222_U29 : ADHALFDL port map( A => mult_222_n50, B => mult_222_n57, CO 
                           => mult_222_n42, S => mult_222_n43);
   mult_222_U28 : ADFULD1 port map( A => mult_222_n64, B => mult_222_n69, CI =>
                           mult_222_n44, CO => mult_222_n40, S => mult_222_n41)
                           ;
   mult_222_U27 : ADFULD1 port map( A => mult_222_n49, B => mult_222_n56, CI =>
                           mult_222_n63, CO => mult_222_n38, S => mult_222_n39)
                           ;
   mult_222_U26 : ADFULD1 port map( A => mult_222_n42, B => mult_222_n68, CI =>
                           mult_222_n39, CO => mult_222_n36, S => mult_222_n37)
                           ;
   mult_222_U24 : ADFULD1 port map( A => mult_222_n55, B => mult_222_n62, CI =>
                           mult_222_n67, CO => mult_222_n32, S => mult_222_n33)
                           ;
   mult_222_U23 : ADFULD1 port map( A => mult_222_n38, B => mult_222_n35, CI =>
                           mult_222_n33, CO => mult_222_n30, S => mult_222_n31)
                           ;
   mult_222_U21 : ADFULD1 port map( A => mult_222_n128, B => mult_222_n61, CI 
                           => mult_222_n54, CO => mult_222_n26, S => 
                           mult_222_n27);
   mult_222_U20 : ADFULD1 port map( A => mult_222_n32, B => mult_222_n29, CI =>
                           mult_222_n27, CO => mult_222_n24, S => mult_222_n25)
                           ;
   mult_222_U18 : ADFULD1 port map( A => mult_222_n126, B => mult_222_n60, CI 
                           => mult_222_n53, CO => mult_222_n20, S => 
                           mult_222_n21);
   mult_222_U17 : ADFULD1 port map( A => mult_222_n26, B => mult_222_n23, CI =>
                           mult_222_n21, CO => mult_222_n18, S => mult_222_n19)
                           ;
   mult_222_U16 : ADFULD1 port map( A => mult_222_n52, B => mult_222_n124, CI 
                           => mult_222_n59, CO => mult_222_n16, S => 
                           mult_222_n17);
   mult_222_U15 : ADFULD1 port map( A => mult_222_n20, B => mult_222_n48, CI =>
                           mult_222_n17, CO => mult_222_n14, S => mult_222_n15)
                           ;
   mult_222_U14 : ADFULD1 port map( A => mult_222_n51, B => mult_222_n47, CI =>
                           mult_222_n16, CO => mult_222_n12, S => mult_222_n13)
                           ;
   mult_222_U13 : ADHALFDL port map( A => mult_222_n71, B => mult_222_n66, CO 
                           => mult_222_n11, S => mult_222_n_1011);
   mult_222_U12 : ADFULD1 port map( A => mult_222_n11, B => mult_222_n58, CI =>
                           mult_222_n45, CO => mult_222_n10, S => 
                           mult_222_n_1010);
   mult_222_U11 : ADFULD1 port map( A => mult_222_n10, B => mult_222_n43, CI =>
                           mult_222_n41, CO => mult_222_n9, S => 
                           mult_222_n_1009);
   mult_222_U10 : ADFULD1 port map( A => mult_222_n37, B => mult_222_n40, CI =>
                           mult_222_n9, CO => mult_222_n8, S => m3_out_6_port);
   mult_222_U9 : ADFULD1 port map( A => mult_222_n31, B => mult_222_n36, CI => 
                           mult_222_n8, CO => mult_222_n7, S => m3_out_7_port);
   mult_222_U8 : ADFULD1 port map( A => mult_222_n25, B => mult_222_n30, CI => 
                           mult_222_n7, CO => mult_222_n6, S => m3_out_8_port);
   mult_222_U7 : ADFULD1 port map( A => mult_222_n19, B => mult_222_n24, CI => 
                           mult_222_n6, CO => mult_222_n5, S => m3_out_9_port);
   mult_222_U6 : ADFULD1 port map( A => mult_222_n15, B => mult_222_n18, CI => 
                           mult_222_n5, CO => mult_222_n4, S => m3_out_10_port)
                           ;
   mult_222_U5 : ADFULD1 port map( A => mult_222_n13, B => mult_222_n14, CI => 
                           mult_222_n4, CO => mult_222_n3, S => m3_out_11_port)
                           ;
   mult_222_U4 : ADFULD1 port map( A => mult_222_n12, B => mult_222_n46, CI => 
                           mult_222_n3, CO => mult_222_n2, S => m3_out_12_port)
                           ;
   mult_221_U201 : EXNOR2D1 port map( A1 => m2_in_r_7_port, A2 => mult_221_n186
                           , Z => mult_221_n197);
   mult_221_U200 : EXOR2D1 port map( A1 => m2_in_r_6_port, A2 => mult_221_n186,
                           Z => mult_221_n211);
   mult_221_U199 : EXNOR2D1 port map( A1 => m2_in_r_7_port, A2 => m2_in_l_5, Z 
                           => mult_221_n204);
   mult_221_U198 : EXOR2D1 port map( A1 => m2_in_r_6_port, A2 => mult_221_n187,
                           Z => mult_221_n203);
   mult_221_U197 : EXNOR2D1 port map( A1 => mult_221_n188, A2 => m3_in_l_0, Z 
                           => mult_221_n86);
   mult_221_U196 : NAN2D1 port map( A1 => mult_221_n212, A2 => mult_221_n86, Z 
                           => mult_221_n37);
   mult_221_U195 : EXNOR2D1 port map( A1 => mult_221_n212, A2 => mult_221_n86, 
                           Z => mult_221_n38);
   mult_221_U194 : NOR2M1D1 port map( A1 => m3_in_l_0, A2 => m2_out_0_port, Z 
                           => mult_221_n60);
   mult_221_U193 : EXNOR2D1 port map( A1 => m2_in_r_5_port, A2 => m3_in_l_0, Z 
                           => mult_221_n210);
   mult_221_U192 : EXNOR2D1 port map( A1 => m2_in_r_4_port, A2 => m3_in_l_0, Z 
                           => mult_221_n209);
   mult_221_U191 : EXNOR2D1 port map( A1 => m2_in_r_3_port, A2 => m3_in_l_0, Z 
                           => mult_221_n208);
   mult_221_U190 : EXNOR2D1 port map( A1 => m2_in_r_2_port, A2 => m3_in_l_0, Z 
                           => mult_221_n207);
   mult_221_U189 : EXNOR2D1 port map( A1 => m2_in_r_1_port, A2 => m3_in_l_0, Z 
                           => mult_221_n206);
   mult_221_U188 : NOR2D1 port map( A1 => mult_221_n205, A2 => mult_221_n194, Z
                           => mult_221_n68);
   mult_221_U187 : EXNOR2D1 port map( A1 => m2_in_r_5_port, A2 => m2_in_l_5, Z 
                           => mult_221_n202);
   mult_221_U186 : EXNOR2D1 port map( A1 => m2_in_r_4_port, A2 => m2_in_l_5, Z 
                           => mult_221_n201);
   mult_221_U185 : EXNOR2D1 port map( A1 => m2_in_r_3_port, A2 => m2_in_l_5, Z 
                           => mult_221_n200);
   mult_221_U184 : EXNOR2D1 port map( A1 => m2_in_r_2_port, A2 => m2_in_l_5, Z 
                           => mult_221_n199);
   mult_221_U183 : EXNOR2D1 port map( A1 => m2_in_r_1_port, A2 => m2_in_l_5, Z 
                           => mult_221_n198);
   mult_221_U182 : NOR2D1 port map( A1 => m2_in_l_5, A2 => mult_221_n194, Z => 
                           mult_221_n76);
   mult_221_U181 : EXNOR2D1 port map( A1 => mult_221_n192, A2 => m3_in_l_0, Z 
                           => mult_221_n87);
   mult_221_U180 : EXNOR2D1 port map( A1 => mult_221_n193, A2 => m3_in_l_0, Z 
                           => mult_221_n88);
   mult_221_U179 : EXOR2D1 port map( A1 => m2_in_r_4_port, A2 => m3_in_l_0, Z 
                           => mult_221_n89);
   mult_221_U178 : EXOR2D1 port map( A1 => m2_in_r_3_port, A2 => m3_in_l_0, Z 
                           => mult_221_n90);
   mult_221_U177 : EXOR2D1 port map( A1 => m2_in_r_2_port, A2 => m3_in_l_0, Z 
                           => mult_221_n91);
   mult_221_U176 : EXOR2D1 port map( A1 => m2_in_r_1_port, A2 => m3_in_l_0, Z 
                           => mult_221_n92);
   mult_221_U175 : EXNOR3D1 port map( A1 => mult_221_n2, A2 => mult_221_n16, A3
                           => mult_221_n196, Z => m2_out_14_port);
   mult_221_U174 : EXOR2D1 port map( A1 => mult_221_n91, A2 => mult_221_n14, Z 
                           => m2_out_2_port);
   mult_221_U173 : EXOR2D1 port map( A1 => mult_221_n75, A2 => mult_221_n53, Z 
                           => mult_221_n50);
   mult_221_U172 : INVD1 port map( A => m2_in_r_7_port, Z => mult_221_n188);
   mult_221_U171 : NOR2D1 port map( A1 => mult_221_n205, A2 => mult_221_n210, Z
                           => mult_221_n63);
   mult_221_U170 : INVD1 port map( A => mult_221_n21, Z => mult_221_n190);
   mult_221_U169 : INVD1 port map( A => m2_in_r_5_port, Z => mult_221_n193);
   mult_221_U168 : INVD1 port map( A => m2_in_r_6_port, Z => mult_221_n192);
   mult_221_U167 : INVD1 port map( A => m2_out_0_port, Z => mult_221_n194);
   mult_221_U166 : NOR2D1 port map( A1 => mult_221_n205, A2 => mult_221_n208, Z
                           => mult_221_n65);
   mult_221_U165 : NOR2D1 port map( A1 => m2_in_l_5, A2 => mult_221_n202, Z => 
                           mult_221_n71);
   mult_221_U164 : NOR2D1 port map( A1 => mult_221_n205, A2 => mult_221_n207, Z
                           => mult_221_n66);
   mult_221_U163 : NOR2D1 port map( A1 => m2_in_l_5, A2 => mult_221_n201, Z => 
                           mult_221_n72);
   mult_221_U162 : NOR2D1 port map( A1 => m2_in_r_4_port, A2 => m3_in_l_0, Z =>
                           mult_221_n79);
   mult_221_U161 : NOR2D1 port map( A1 => m2_in_l_5, A2 => mult_221_n198, Z => 
                           mult_221_n75);
   mult_221_U160 : NOR2D1 port map( A1 => m2_in_r_2_port, A2 => m3_in_l_0, Z =>
                           mult_221_n81);
   mult_221_U159 : NOR2D1 port map( A1 => mult_221_n205, A2 => mult_221_n206, Z
                           => mult_221_n67);
   mult_221_U158 : NOR3D1 port map( A1 => mult_221_n205, A2 => mult_221_n186, 
                           A3 => m2_out_0_port, Z => mult_221_n57);
   mult_221_U157 : NOR2D1 port map( A1 => m2_in_l_5, A2 => mult_221_n200, Z => 
                           mult_221_n73);
   mult_221_U156 : NOR2D1 port map( A1 => m2_in_r_1_port, A2 => m3_in_l_0, Z =>
                           mult_221_n82);
   mult_221_U155 : NOR2D1 port map( A1 => m2_in_r_3_port, A2 => m3_in_l_0, Z =>
                           mult_221_n80);
   mult_221_U154 : NOR2D1 port map( A1 => m2_in_l_5, A2 => mult_221_n199, Z => 
                           mult_221_n74);
   mult_221_U153 : NOR2D1 port map( A1 => m2_out_0_port, A2 => m3_in_l_0, Z => 
                           mult_221_n83);
   mult_221_U152 : NAN2D1 port map( A1 => mult_221_n195, A2 => mult_221_n197, Z
                           => mult_221_n196);
   mult_221_U151 : NAN2D1 port map( A1 => mult_221_n195, A2 => mult_221_n197, Z
                           => mult_221_n16);
   mult_221_U150 : INVD1 port map( A => mult_221_n204, Z => mult_221_n189);
   mult_221_U149 : NOR2D1 port map( A1 => mult_221_n205, A2 => mult_221_n211, Z
                           => mult_221_n62);
   mult_221_U148 : NAN2D1 port map( A1 => mult_221_n187, A2 => mult_221_n189, Z
                           => mult_221_n69);
   mult_221_U147 : NOR2D1 port map( A1 => m2_in_l_5, A2 => mult_221_n204, Z => 
                           mult_221_n21);
   mult_221_U146 : NOR2D1 port map( A1 => mult_221_n205, A2 => mult_221_n209, Z
                           => mult_221_n64);
   mult_221_U145 : INVD1 port map( A => mult_221_n32, Z => mult_221_n191);
   mult_221_U144 : NOR2D1 port map( A1 => m2_in_l_5, A2 => mult_221_n203, Z => 
                           mult_221_n70);
   mult_221_U143 : NAN2D1 port map( A1 => mult_221_n186, A2 => mult_221_n188, Z
                           => mult_221_n77);
   mult_221_U142 : NAN2D1 port map( A1 => mult_221_n192, A2 => mult_221_n186, Z
                           => mult_221_n32);
   mult_221_U141 : NAN2D1 port map( A1 => mult_221_n193, A2 => mult_221_n186, Z
                           => mult_221_n212);
   mult_221_U140 : INVD1 port map( A => m2_in_l_5, Z => mult_221_n187);
   mult_221_U139 : EXOR2D1 port map( A1 => m3_in_l_0, A2 => mult_221_n187, Z =>
                           mult_221_n205);
   mult_221_U138 : INVD1 port map( A => m3_in_l_0, Z => mult_221_n186);
   mult_221_U137 : AND2D1 port map( A1 => mult_221_n53, A2 => mult_221_n75, Z 
                           => mult_221_n185);
   mult_221_U136 : INVD1 port map( A => mult_221_n205, Z => mult_221_n195);
   mult_221_U135 : AND2D1 port map( A1 => mult_221_n14, A2 => mult_221_n91, Z 
                           => mult_221_n184);
   mult_221_U37 : ADHALFDL port map( A => mult_221_n186, B => mult_221_n90, CO 
                           => mult_221_n55, S => mult_221_n56);
   mult_221_U36 : ADFULD1 port map( A => mult_221_n89, B => mult_221_n76, CI =>
                           mult_221_n82, CO => mult_221_n53, S => mult_221_n54)
                           ;
   mult_221_U35 : ADHALFDL port map( A => mult_221_n81, B => mult_221_n88, CO 
                           => mult_221_n51, S => mult_221_n52);
   mult_221_U33 : ADFULD1 port map( A => mult_221_n68, B => mult_221_n87, CI =>
                           mult_221_n80, CO => mult_221_n47, S => mult_221_n48)
                           ;
   mult_221_U32 : ADFULD1 port map( A => mult_221_n51, B => mult_221_n74, CI =>
                           mult_221_n48, CO => mult_221_n45, S => mult_221_n46)
                           ;
   mult_221_U31 : ADHALFDL port map( A => mult_221_n79, B => mult_221_n86, CO 
                           => mult_221_n43, S => mult_221_n44);
   mult_221_U30 : ADFULD1 port map( A => mult_221_n67, B => mult_221_n73, CI =>
                           mult_221_n57, CO => mult_221_n41, S => mult_221_n42)
                           ;
   mult_221_U29 : ADFULD1 port map( A => mult_221_n44, B => mult_221_n47, CI =>
                           mult_221_n42, CO => mult_221_n39, S => mult_221_n40)
                           ;
   mult_221_U26 : ADFULD1 port map( A => mult_221_n66, B => mult_221_n72, CI =>
                           mult_221_n43, CO => mult_221_n35, S => mult_221_n36)
                           ;
   mult_221_U25 : ADFULD1 port map( A => mult_221_n41, B => mult_221_n38, CI =>
                           mult_221_n36, CO => mult_221_n33, S => mult_221_n34)
                           ;
   mult_221_U23 : ADFULD1 port map( A => mult_221_n65, B => mult_221_n71, CI =>
                           mult_221_n32, CO => mult_221_n29, S => mult_221_n30)
                           ;
   mult_221_U22 : ADFULD1 port map( A => mult_221_n35, B => mult_221_n37, CI =>
                           mult_221_n30, CO => mult_221_n27, S => mult_221_n28)
                           ;
   mult_221_U21 : ADFULD1 port map( A => mult_221_n70, B => mult_221_n191, CI 
                           => mult_221_n64, CO => mult_221_n25, S => 
                           mult_221_n26);
   mult_221_U20 : ADFULD1 port map( A => mult_221_n29, B => mult_221_n77, CI =>
                           mult_221_n26, CO => mult_221_n23, S => mult_221_n24)
                           ;
   mult_221_U18 : ADFULD1 port map( A => mult_221_n190, B => mult_221_n63, CI 
                           => mult_221_n25, CO => mult_221_n19, S => 
                           mult_221_n20);
   mult_221_U17 : ADFULD1 port map( A => mult_221_n62, B => mult_221_n21, CI =>
                           mult_221_n69, CO => mult_221_n17, S => mult_221_n18)
                           ;
   mult_221_U15 : ADHALFDL port map( A => mult_221_n92, B => mult_221_n60, CO 
                           => mult_221_n14, S => m2_out_1_port);
   mult_221_U13 : ADFULD1 port map( A => mult_221_n56, B => mult_221_n83, CI =>
                           mult_221_n184, CO => mult_221_n12, S => 
                           m2_out_3_port);
   mult_221_U12 : ADFULD1 port map( A => mult_221_n54, B => mult_221_n55, CI =>
                           mult_221_n12, CO => mult_221_n11, S => m2_out_4_port
                           );
   mult_221_U11 : ADFULD1 port map( A => mult_221_n50, B => mult_221_n52, CI =>
                           mult_221_n11, CO => mult_221_n10, S => m2_out_5_port
                           );
   mult_221_U10 : ADFULD1 port map( A => mult_221_n46, B => mult_221_n185, CI 
                           => mult_221_n10, CO => mult_221_n9, S => 
                           m2_out_6_port);
   mult_221_U9 : ADFULD1 port map( A => mult_221_n40, B => mult_221_n45, CI => 
                           mult_221_n9, CO => mult_221_n8, S => m2_out_7_port);
   mult_221_U8 : ADFULD1 port map( A => mult_221_n34, B => mult_221_n39, CI => 
                           mult_221_n8, CO => mult_221_n7, S => m2_out_8_port);
   mult_221_U7 : ADFULD1 port map( A => mult_221_n28, B => mult_221_n33, CI => 
                           mult_221_n7, CO => mult_221_n6, S => m2_out_9_port);
   mult_221_U6 : ADFULD1 port map( A => mult_221_n24, B => mult_221_n27, CI => 
                           mult_221_n6, CO => mult_221_n5, S => m2_out_10_port)
                           ;
   mult_221_U5 : ADFULD1 port map( A => mult_221_n20, B => mult_221_n23, CI => 
                           mult_221_n5, CO => mult_221_n4, S => m2_out_11_port)
                           ;
   mult_221_U4 : ADFULD1 port map( A => mult_221_n19, B => mult_221_n18, CI => 
                           mult_221_n4, CO => mult_221_n3, S => m2_out_12_port)
                           ;
   mult_221_U3 : ADFULD1 port map( A => mult_221_n17, B => mult_221_n16, CI => 
                           mult_221_n3, CO => mult_221_n2, S => m2_out_13_port)
                           ;
   mult_220_U159 : MUX2DL port map( A0 => mult_220_n177, A1 => mult_220_n176, 
                           SL => m3_in_l_0, Z => mult_220_n106);
   mult_220_U158 : MUX2DL port map( A0 => mult_220_n179, A1 => mult_220_n177, 
                           SL => m3_in_l_0, Z => mult_220_n107);
   mult_220_U157 : MUX2DL port map( A0 => mult_220_n180, A1 => mult_220_n179, 
                           SL => m3_in_l_0, Z => mult_220_n108);
   mult_220_U156 : MUX2DL port map( A0 => mult_220_n181, A1 => mult_220_n180, 
                           SL => m3_in_l_0, Z => mult_220_n109);
   mult_220_U155 : MUX2DL port map( A0 => mult_220_n182, A1 => mult_220_n181, 
                           SL => m3_in_l_0, Z => mult_220_n110);
   mult_220_U154 : MUX2DL port map( A0 => mult_220_n183, A1 => mult_220_n182, 
                           SL => m3_in_l_0, Z => mult_220_n111);
   mult_220_U153 : MUX2DL port map( A0 => mult_220_n185, A1 => mult_220_n183, 
                           SL => m3_in_l_0, Z => mult_220_n112);
   mult_220_U152 : NAN2D1 port map( A1 => m3_in_l_0, A2 => m1_in_r_0_port, Z =>
                           mult_220_n15);
   mult_220_U151 : MUX2DL port map( A0 => mult_220_n177, A1 => mult_220_n176, 
                           SL => m3_in_l_0, Z => mult_220_n55);
   mult_220_U150 : MUX2DL port map( A0 => mult_220_n179, A1 => mult_220_n177, 
                           SL => m3_in_l_0, Z => mult_220_n56);
   mult_220_U149 : MUX2DL port map( A0 => mult_220_n180, A1 => mult_220_n179, 
                           SL => m3_in_l_0, Z => mult_220_n57);
   mult_220_U148 : MUX2DL port map( A0 => mult_220_n181, A1 => mult_220_n180, 
                           SL => m3_in_l_0, Z => mult_220_n58);
   mult_220_U147 : MUX2DL port map( A0 => mult_220_n182, A1 => mult_220_n181, 
                           SL => m3_in_l_0, Z => mult_220_n59);
   mult_220_U146 : MUX2DL port map( A0 => mult_220_n183, A1 => mult_220_n182, 
                           SL => m3_in_l_0, Z => mult_220_n60);
   mult_220_U145 : MUX2DL port map( A0 => mult_220_n185, A1 => mult_220_n183, 
                           SL => m3_in_l_0, Z => mult_220_n61);
   mult_220_U144 : NAN2D1 port map( A1 => m3_in_l_0, A2 => m1_in_r_0_port, Z =>
                           mult_220_n62);
   mult_220_U143 : NAN2M1D1 port map( A1 => mult_220_n174, A2 => m1_in_r_7_port
                           , Z => mult_220_n88);
   mult_220_U142 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => m1_in_r_7_port, Z 
                           => mult_220_n97);
   mult_220_U141 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n176, Z => mult_220_n187);
   mult_220_U140 : EXNOR3D1 port map( A1 => mult_220_n2, A2 => mult_220_n16, A3
                           => mult_220_n187, Z => m1_out_14_port);
   mult_220_U139 : TIEHI port map( Z => mult_220_n186);
   mult_220_U138 : INVD1 port map( A => m1_in_r_7_port, Z => mult_220_n176);
   mult_220_U137 : INVD1 port map( A => m1_in_r_6_port, Z => mult_220_n177);
   mult_220_U136 : INVD1 port map( A => m1_in_r_5_port, Z => mult_220_n179);
   mult_220_U135 : INVD1 port map( A => m1_in_r_4_port, Z => mult_220_n180);
   mult_220_U134 : INVD1 port map( A => m1_in_r_3_port, Z => mult_220_n181);
   mult_220_U133 : INVD1 port map( A => m1_in_r_2_port, Z => mult_220_n182);
   mult_220_U132 : INVD1 port map( A => m1_in_r_1_port, Z => mult_220_n183);
   mult_220_U131 : INVD1 port map( A => m1_in_r_0_port, Z => mult_220_n185);
   mult_220_U130 : INVD1 port map( A => mult_220_n15, Z => m1_out_0_port);
   mult_220_U129 : INVD1 port map( A => mult_220_n22, Z => mult_220_n178);
   mult_220_U128 : INVD1 port map( A => mult_220_n16, Z => mult_220_n175);
   mult_220_U127 : NAN2D1 port map( A1 => m3_in_l_0, A2 => mult_220_n174, Z => 
                           mult_220_n126);
   mult_220_U126 : INVD1 port map( A => m2_in_l_5, Z => mult_220_n174);
   mult_220_U88 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => mult_220_n185, Z =>
                           mult_220_n105);
   mult_220_U86 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => mult_220_n183, Z =>
                           mult_220_n104);
   mult_220_U84 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => mult_220_n182, Z =>
                           mult_220_n103);
   mult_220_U82 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => mult_220_n181, Z =>
                           mult_220_n102);
   mult_220_U80 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => mult_220_n180, Z =>
                           mult_220_n101);
   mult_220_U78 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => mult_220_n179, Z =>
                           mult_220_n100);
   mult_220_U76 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => mult_220_n177, Z =>
                           mult_220_n99);
   mult_220_U74 : EXNOR2D1 port map( A1 => m2_in_l_5, A2 => mult_220_n176, Z =>
                           mult_220_n98);
   mult_220_U70 : NOR2D1 port map( A1 => mult_220_n186, A2 => mult_220_n174, Z 
                           => mult_220_n96);
   mult_220_U68 : NOR2D1 port map( A1 => mult_220_n185, A2 => mult_220_n174, Z 
                           => mult_220_n95);
   mult_220_U66 : NOR2D1 port map( A1 => mult_220_n183, A2 => mult_220_n174, Z 
                           => mult_220_n94);
   mult_220_U64 : NOR2D1 port map( A1 => mult_220_n182, A2 => mult_220_n174, Z 
                           => mult_220_n93);
   mult_220_U62 : NOR2D1 port map( A1 => mult_220_n181, A2 => mult_220_n174, Z 
                           => mult_220_n92);
   mult_220_U60 : NOR2D1 port map( A1 => mult_220_n180, A2 => mult_220_n174, Z 
                           => mult_220_n91);
   mult_220_U58 : NOR2D1 port map( A1 => mult_220_n179, A2 => mult_220_n174, Z 
                           => mult_220_n90);
   mult_220_U56 : NOR2D1 port map( A1 => mult_220_n177, A2 => mult_220_n174, Z 
                           => mult_220_n89);
   mult_220_U53 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n62, Z => mult_220_n87);
   mult_220_U51 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n61, Z => mult_220_n86);
   mult_220_U49 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n60, Z => mult_220_n85);
   mult_220_U47 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n59, Z => mult_220_n84);
   mult_220_U45 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n58, Z => mult_220_n83);
   mult_220_U43 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n57, Z => mult_220_n22);
   mult_220_U41 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n56, Z => mult_220_n82);
   mult_220_U39 : MUXB2DL port map( A0 => mult_220_n126, A1 => mult_220_n174, 
                           SL => mult_220_n55, Z => mult_220_n16);
   mult_220_U36 : ADHALFDL port map( A => mult_220_n111, B => m2_in_l_5, CO => 
                           mult_220_n53, S => mult_220_n54);
   mult_220_U35 : ADHALFDL port map( A => mult_220_n104, B => mult_220_n110, CO
                           => mult_220_n51, S => mult_220_n52);
   mult_220_U34 : ADFULD1 port map( A => mult_220_n103, B => mult_220_n109, CI 
                           => mult_220_n96, CO => mult_220_n49, S => 
                           mult_220_n50);
   mult_220_U33 : ADFULD1 port map( A => mult_220_n102, B => mult_220_n108, CI 
                           => mult_220_n95, CO => mult_220_n47, S => 
                           mult_220_n48);
   mult_220_U32 : ADFULD1 port map( A => m2_in_l_5, B => mult_220_n107, CI => 
                           mult_220_n101, CO => mult_220_n45, S => mult_220_n46
                           );
   mult_220_U31 : ADFULD1 port map( A => mult_220_n94, B => mult_220_n87, CI =>
                           mult_220_n46, CO => mult_220_n43, S => mult_220_n44)
                           ;
   mult_220_U30 : ADFULD1 port map( A => mult_220_n100, B => mult_220_n106, CI 
                           => mult_220_n86, CO => mult_220_n41, S => 
                           mult_220_n42);
   mult_220_U29 : ADFULD1 port map( A => mult_220_n45, B => mult_220_n93, CI =>
                           mult_220_n42, CO => mult_220_n39, S => mult_220_n40)
                           ;
   mult_220_U27 : ADFULD1 port map( A => mult_220_n99, B => mult_220_n176, CI 
                           => mult_220_n85, CO => mult_220_n36, S => 
                           mult_220_n37);
   mult_220_U26 : ADFULD1 port map( A => mult_220_n41, B => mult_220_n92, CI =>
                           mult_220_n37, CO => mult_220_n34, S => mult_220_n35)
                           ;
   mult_220_U24 : ADFULD1 port map( A => mult_220_n98, B => mult_220_n176, CI 
                           => mult_220_n84, CO => mult_220_n30, S => 
                           mult_220_n31);
   mult_220_U23 : ADFULD1 port map( A => mult_220_n36, B => mult_220_n91, CI =>
                           mult_220_n31, CO => mult_220_n28, S => mult_220_n29)
                           ;
   mult_220_U22 : ADFULD1 port map( A => mult_220_n97, B => m1_in_r_7_port, CI 
                           => mult_220_n83, CO => mult_220_n26, S => 
                           mult_220_n27);
   mult_220_U21 : ADFULD1 port map( A => mult_220_n30, B => mult_220_n90, CI =>
                           mult_220_n27, CO => mult_220_n24, S => mult_220_n25)
                           ;
   mult_220_U19 : ADFULD1 port map( A => mult_220_n178, B => mult_220_n89, CI 
                           => mult_220_n26, CO => mult_220_n20, S => 
                           mult_220_n21);
   mult_220_U18 : ADFULD1 port map( A => mult_220_n82, B => mult_220_n88, CI =>
                           mult_220_n22, CO => mult_220_n18, S => mult_220_n19)
                           ;
   mult_220_U15 : ADHALFDL port map( A => mult_220_n112, B => mult_220_n15, CO 
                           => mult_220_n14, S => m1_out_1_port);
   mult_220_U14 : ADFULD1 port map( A => mult_220_n14, B => mult_220_n105, CI 
                           => mult_220_n54, CO => mult_220_n13, S => 
                           m1_out_2_port);
   mult_220_U13 : ADFULD1 port map( A => mult_220_n52, B => mult_220_n53, CI =>
                           mult_220_n13, CO => mult_220_n12, S => m1_out_3_port
                           );
   mult_220_U12 : ADFULD1 port map( A => mult_220_n50, B => mult_220_n51, CI =>
                           mult_220_n12, CO => mult_220_n11, S => m1_out_4_port
                           );
   mult_220_U11 : ADFULD1 port map( A => mult_220_n48, B => mult_220_n49, CI =>
                           mult_220_n11, CO => mult_220_n10, S => m1_out_5_port
                           );
   mult_220_U10 : ADFULD1 port map( A => mult_220_n44, B => mult_220_n47, CI =>
                           mult_220_n10, CO => mult_220_n9, S => m1_out_6_port)
                           ;
   mult_220_U9 : ADFULD1 port map( A => mult_220_n40, B => mult_220_n43, CI => 
                           mult_220_n9, CO => mult_220_n8, S => m1_out_7_port);
   mult_220_U8 : ADFULD1 port map( A => mult_220_n35, B => mult_220_n39, CI => 
                           mult_220_n8, CO => mult_220_n7, S => m1_out_8_port);
   mult_220_U7 : ADFULD1 port map( A => mult_220_n29, B => mult_220_n34, CI => 
                           mult_220_n7, CO => mult_220_n6, S => m1_out_9_port);
   mult_220_U6 : ADFULD1 port map( A => mult_220_n25, B => mult_220_n28, CI => 
                           mult_220_n6, CO => mult_220_n5, S => m1_out_10_port)
                           ;
   mult_220_U5 : ADFULD1 port map( A => mult_220_n21, B => mult_220_n24, CI => 
                           mult_220_n5, CO => mult_220_n4, S => m1_out_11_port)
                           ;
   mult_220_U4 : ADFULD1 port map( A => mult_220_n20, B => mult_220_n19, CI => 
                           mult_220_n4, CO => mult_220_n3, S => m1_out_12_port)
                           ;
   mult_220_U3 : ADFULD1 port map( A => mult_220_n18, B => mult_220_n175, CI =>
                           mult_220_n3, CO => mult_220_n2, S => m1_out_13_port)
                           ;

end flat_rtl_none_10;
