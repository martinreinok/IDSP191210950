
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_sec_nov_std is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_sec_nov_std;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_sec_nov_std.all;

architecture flat_rtl_none_10 of sec_nov_std is

   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AO21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3M1D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component NAN4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   signal sec_nov_inst_n_1017, sec_nov_inst_n_1016, sec_nov_inst_n_1015, 
      sec_nov_inst_n_1014, sec_nov_inst_n_1013, sec_nov_inst_n_1012, 
      sec_nov_inst_n_1011, sec_nov_inst_n_1010, sec_nov_inst_n85, 
      sec_nov_inst_n58, sec_nov_inst_n51, sec_nov_inst_n50, sec_nov_inst_n49, 
      sec_nov_inst_n48, sec_nov_inst_n47, sec_nov_inst_n46, sec_nov_inst_n45, 
      sec_nov_inst_n44, sec_nov_inst_n43, sec_nov_inst_n42, sec_nov_inst_n41, 
      sec_nov_inst_n40, sec_nov_inst_n39, sec_nov_inst_n38, sec_nov_inst_n37, 
      sec_nov_inst_n36, sec_nov_inst_n35, sec_nov_inst_n34, sec_nov_inst_n33, 
      sec_nov_inst_n32, sec_nov_inst_n31, sec_nov_inst_n30, sec_nov_inst_n29, 
      sec_nov_inst_n28, sec_nov_inst_n27, sec_nov_inst_n26, sec_nov_inst_n25, 
      sec_nov_inst_n24, sec_nov_inst_n23, sec_nov_inst_n22, sec_nov_inst_n21, 
      sec_nov_inst_n20, sec_nov_inst_n19, sec_nov_inst_n18, sec_nov_inst_n17, 
      sec_nov_inst_n16, sec_nov_inst_n15, sec_nov_inst_n14, sec_nov_inst_n13, 
      sec_nov_inst_n12, sec_nov_inst_n11, sec_nov_inst_n10, sec_nov_inst_n9, 
      sec_nov_inst_n8, sec_nov_inst_n6, sec_nov_inst_n5, sec_nov_inst_n4, 
      sec_nov_inst_n3, sec_nov_inst_n2, sec_nov_inst_n1, 
      sec_nov_inst_add_416_C239_rn_carry_7_port, 
      sec_nov_inst_add_416_C239_rn_carry_6_port, 
      sec_nov_inst_add_416_C239_rn_carry_5_port, 
      sec_nov_inst_add_416_C239_rn_carry_4_port, 
      sec_nov_inst_add_416_C239_rn_carry_3_port, 
      sec_nov_inst_add_416_C239_rn_carry_2_port, 
      sec_nov_inst_add_416_C239_rn_carry_1_port, sec_nov_inst_n84, 
      sec_nov_inst_n83, sec_nov_inst_n82, sec_nov_inst_n81, sec_nov_inst_n80, 
      sec_nov_inst_n79, sec_nov_inst_n78, sec_nov_inst_n77, sec_nov_inst_n76, 
      sec_nov_inst_n75, sec_nov_inst_n74, sec_nov_inst_n73, sec_nov_inst_n72, 
      sec_nov_inst_n71, sec_nov_inst_n70, sec_nov_inst_n69, sec_nov_inst_n68, 
      sec_nov_inst_n67, sec_nov_inst_n66, sec_nov_inst_n65, sec_nov_inst_n64, 
      sec_nov_inst_n63, sec_nov_inst_n62, sec_nov_inst_n61, sec_nov_inst_n60, 
      sec_nov_inst_n59, sec_nov_inst_n57, sec_nov_inst_n56, sec_nov_inst_n55, 
      sec_nov_inst_n54, sec_nov_inst_n53, sec_nov_inst_n52, sec_nov_inst_n7, 
      sec_nov_inst_N131, sec_nov_inst_N130, sec_nov_inst_N129, 
      sec_nov_inst_N128, sec_nov_inst_N127, sec_nov_inst_N126, 
      sec_nov_inst_N125, sec_nov_inst_N124, sec_nov_inst_N123, 
      sec_nov_inst_state_0_port, sec_nov_inst_state_1_port, 
      sec_nov_inst_state_2_port, sec_nov_inst_state_3_port, 
      sec_nov_inst_a_out_0_port, sec_nov_inst_a_out_1_port, 
      sec_nov_inst_a_out_2_port, sec_nov_inst_a_out_3_port, 
      sec_nov_inst_a_out_4_port, sec_nov_inst_a_out_5_port, 
      sec_nov_inst_a_out_6_port, sec_nov_inst_a_out_7_port, 
      sec_nov_inst_a_in_r_0_port, sec_nov_inst_a_in_r_1_port, 
      sec_nov_inst_a_in_r_2_port, sec_nov_inst_a_in_r_3_port, 
      sec_nov_inst_a_in_r_4_port, sec_nov_inst_a_in_r_5_port, 
      sec_nov_inst_a_in_r_6_port, sec_nov_inst_a_in_r_7_port, 
      sec_nov_inst_a_in_r_8_port, sec_nov_inst_a_in_r_9_port, 
      sec_nov_inst_a_in_r_10_port, sec_nov_inst_a_in_r_11_port, 
      sec_nov_inst_a_in_r_12_port, sec_nov_inst_a_in_r_13_port, 
      sec_nov_inst_a_in_r_14_port, sec_nov_inst_a_in_l_0_port, 
      sec_nov_inst_a_in_l_1_port, sec_nov_inst_a_in_l_2_port, 
      sec_nov_inst_a_in_l_3_port, sec_nov_inst_a_in_l_4_port, 
      sec_nov_inst_a_in_l_5_port, sec_nov_inst_a_in_l_6_port, 
      sec_nov_inst_a_in_l_7_port, sec_nov_inst_a_in_l_8_port, 
      sec_nov_inst_a_in_l_9_port, sec_nov_inst_a_in_l_10_port, 
      sec_nov_inst_a_in_l_11_port, sec_nov_inst_a_in_l_12_port, 
      sec_nov_inst_a_in_l_13_port, sec_nov_inst_a_in_l_14_port, 
      sec_nov_inst_m_out_0_port, sec_nov_inst_m_out_1_port, 
      sec_nov_inst_m_out_2_port, sec_nov_inst_m_out_3_port, 
      sec_nov_inst_m_out_4_port, sec_nov_inst_m_out_5_port, 
      sec_nov_inst_m_out_6_port, sec_nov_inst_m_out_7_port, 
      sec_nov_inst_m_out_8_port, sec_nov_inst_m_out_9_port, 
      sec_nov_inst_m_out_10_port, sec_nov_inst_m_out_11_port, 
      sec_nov_inst_m_out_12_port, sec_nov_inst_m_out_13_port, 
      sec_nov_inst_m_out_14_port, sec_nov_inst_m_in_r_0_port, 
      sec_nov_inst_m_in_r_1_port, sec_nov_inst_m_in_r_2_port, 
      sec_nov_inst_m_in_r_3_port, sec_nov_inst_m_in_r_4_port, 
      sec_nov_inst_m_in_r_5_port, sec_nov_inst_m_in_r_6_port, 
      sec_nov_inst_m_in_r_7_port, sec_nov_inst_m_in_l_0_port, 
      sec_nov_inst_m_in_l_1_port, sec_nov_inst_m_in_l_2_port, 
      sec_nov_inst_m_in_l_3_port, sec_nov_inst_m_in_l_4_port, 
      sec_nov_inst_m_in_l_5_port, sec_nov_inst_m_in_l_6_port, 
      sec_nov_inst_m_in_l_7_port, sec_nov_inst_arx_state_reg_0_port, 
      sec_nov_inst_arx_state_reg_1_port, sec_nov_inst_arx_state_reg_2_port, 
      sec_nov_inst_arx_state_reg_3_port, sec_nov_inst_arx_d2_reg_0_port, 
      sec_nov_inst_arx_d2_reg_1_port, sec_nov_inst_arx_d2_reg_2_port, 
      sec_nov_inst_arx_d2_reg_3_port, sec_nov_inst_arx_d2_reg_4_port, 
      sec_nov_inst_arx_d2_reg_5_port, sec_nov_inst_arx_d2_reg_6_port, 
      sec_nov_inst_arx_d2_reg_7_port, sec_nov_inst_arx_d1_reg_0_port, 
      sec_nov_inst_arx_d1_reg_1_port, sec_nov_inst_arx_d1_reg_2_port, 
      sec_nov_inst_arx_d1_reg_3_port, sec_nov_inst_arx_d1_reg_4_port, 
      sec_nov_inst_arx_d1_reg_5_port, sec_nov_inst_arx_d1_reg_6_port, 
      sec_nov_inst_arx_d1_reg_7_port, sec_nov_inst_arx_d0_reg_0_port, 
      sec_nov_inst_arx_d0_reg_1_port, sec_nov_inst_arx_d0_reg_2_port, 
      sec_nov_inst_arx_d0_reg_3_port, sec_nov_inst_arx_d0_reg_4_port, 
      sec_nov_inst_arx_d0_reg_5_port, sec_nov_inst_arx_d0_reg_6_port, 
      sec_nov_inst_arx_d0_reg_7_port, sec_nov_inst_arx_r4_reg_0_port, 
      sec_nov_inst_arx_r4_reg_1_port, sec_nov_inst_arx_r4_reg_2_port, 
      sec_nov_inst_arx_r4_reg_3_port, sec_nov_inst_arx_r4_reg_4_port, 
      sec_nov_inst_arx_r4_reg_5_port, sec_nov_inst_arx_r4_reg_6_port, 
      sec_nov_inst_arx_r4_reg_7_port, sec_nov_inst_arx_r3_reg_0_port, 
      sec_nov_inst_arx_r3_reg_1_port, sec_nov_inst_arx_r3_reg_2_port, 
      sec_nov_inst_arx_r3_reg_3_port, sec_nov_inst_arx_r3_reg_4_port, 
      sec_nov_inst_arx_r3_reg_5_port, sec_nov_inst_arx_r3_reg_6_port, 
      sec_nov_inst_arx_r3_reg_7_port, sec_nov_inst_arx_r3_reg_8_port, 
      sec_nov_inst_arx_r3_reg_9_port, sec_nov_inst_arx_r3_reg_10_port, 
      sec_nov_inst_arx_r3_reg_11_port, sec_nov_inst_arx_r3_reg_12_port, 
      sec_nov_inst_arx_r3_reg_13_port, sec_nov_inst_arx_r3_reg_14_port, 
      sec_nov_inst_arx_r2_reg_0_port, sec_nov_inst_arx_r2_reg_1_port, 
      sec_nov_inst_arx_r2_reg_2_port, sec_nov_inst_arx_r2_reg_3_port, 
      sec_nov_inst_arx_r2_reg_4_port, sec_nov_inst_arx_r2_reg_5_port, 
      sec_nov_inst_arx_r2_reg_6_port, sec_nov_inst_arx_r2_reg_7_port, 
      sec_nov_inst_arx_r2_reg_8_port, sec_nov_inst_arx_r2_reg_9_port, 
      sec_nov_inst_arx_r2_reg_10_port, sec_nov_inst_arx_r2_reg_11_port, 
      sec_nov_inst_arx_r2_reg_12_port, sec_nov_inst_arx_r2_reg_13_port, 
      sec_nov_inst_arx_r2_reg_14_port, sec_nov_inst_arx_r1_reg_0_port, 
      sec_nov_inst_arx_r1_reg_1_port, sec_nov_inst_arx_r1_reg_2_port, 
      sec_nov_inst_arx_r1_reg_3_port, sec_nov_inst_arx_r1_reg_4_port, 
      sec_nov_inst_arx_r1_reg_5_port, sec_nov_inst_arx_r1_reg_6_port, 
      sec_nov_inst_arx_r1_reg_7_port, sec_nov_inst_arx_i1_reg_0_port, 
      sec_nov_inst_arx_i1_reg_1_port, sec_nov_inst_arx_i1_reg_2_port, 
      sec_nov_inst_arx_i1_reg_3_port, sec_nov_inst_arx_i1_reg_4_port, 
      sec_nov_inst_arx_i1_reg_5_port, sec_nov_inst_arx_i1_reg_6_port, 
      sec_nov_inst_arx_i1_reg_7_port, sec_nov_inst_add_239_n_1009, 
      sec_nov_inst_add_239_n9, sec_nov_inst_add_239_n8, sec_nov_inst_add_239_n7
      , sec_nov_inst_add_239_n6, sec_nov_inst_add_239_n5, 
      sec_nov_inst_add_239_n4, sec_nov_inst_add_239_n3, sec_nov_inst_add_239_n2
      , sec_nov_inst_add_239_n1, sec_nov_inst_add_239_carry_6_port, 
      sec_nov_inst_add_239_carry_7_port, sec_nov_inst_add_239_carry_8_port, 
      sec_nov_inst_add_239_carry_9_port, sec_nov_inst_add_239_carry_10_port, 
      sec_nov_inst_add_239_carry_11_port, sec_nov_inst_add_239_carry_12_port, 
      sec_nov_inst_add_239_carry_13_port, sec_nov_inst_add_239_carry_14_port, 
      sec_nov_inst_mult_238_n247, sec_nov_inst_mult_238_n246, 
      sec_nov_inst_mult_238_n245, sec_nov_inst_mult_238_n244, 
      sec_nov_inst_mult_238_n243, sec_nov_inst_mult_238_n242, 
      sec_nov_inst_mult_238_n241, sec_nov_inst_mult_238_n240, 
      sec_nov_inst_mult_238_n239, sec_nov_inst_mult_238_n238, 
      sec_nov_inst_mult_238_n237, sec_nov_inst_mult_238_n236, 
      sec_nov_inst_mult_238_n235, sec_nov_inst_mult_238_n234, 
      sec_nov_inst_mult_238_n233, sec_nov_inst_mult_238_n232, 
      sec_nov_inst_mult_238_n231, sec_nov_inst_mult_238_n230, 
      sec_nov_inst_mult_238_n229, sec_nov_inst_mult_238_n228, 
      sec_nov_inst_mult_238_n227, sec_nov_inst_mult_238_n226, 
      sec_nov_inst_mult_238_n225, sec_nov_inst_mult_238_n224, 
      sec_nov_inst_mult_238_n223, sec_nov_inst_mult_238_n222, 
      sec_nov_inst_mult_238_n221, sec_nov_inst_mult_238_n220, 
      sec_nov_inst_mult_238_n219, sec_nov_inst_mult_238_n218, 
      sec_nov_inst_mult_238_n217, sec_nov_inst_mult_238_n216, 
      sec_nov_inst_mult_238_n215, sec_nov_inst_mult_238_n214, 
      sec_nov_inst_mult_238_n213, sec_nov_inst_mult_238_n212, 
      sec_nov_inst_mult_238_n211, sec_nov_inst_mult_238_n210, 
      sec_nov_inst_mult_238_n209, sec_nov_inst_mult_238_n208, 
      sec_nov_inst_mult_238_n207, sec_nov_inst_mult_238_n206, 
      sec_nov_inst_mult_238_n205, sec_nov_inst_mult_238_n204, 
      sec_nov_inst_mult_238_n203, sec_nov_inst_mult_238_n202, 
      sec_nov_inst_mult_238_n201, sec_nov_inst_mult_238_n200, 
      sec_nov_inst_mult_238_n199, sec_nov_inst_mult_238_n198, 
      sec_nov_inst_mult_238_n197, sec_nov_inst_mult_238_n196, 
      sec_nov_inst_mult_238_n195, sec_nov_inst_mult_238_n194, 
      sec_nov_inst_mult_238_n92, sec_nov_inst_mult_238_n91, 
      sec_nov_inst_mult_238_n90, sec_nov_inst_mult_238_n89, 
      sec_nov_inst_mult_238_n88, sec_nov_inst_mult_238_n87, 
      sec_nov_inst_mult_238_n86, sec_nov_inst_mult_238_n85, 
      sec_nov_inst_mult_238_n84, sec_nov_inst_mult_238_n83, 
      sec_nov_inst_mult_238_n82, sec_nov_inst_mult_238_n81, 
      sec_nov_inst_mult_238_n80, sec_nov_inst_mult_238_n79, 
      sec_nov_inst_mult_238_n77, sec_nov_inst_mult_238_n76, 
      sec_nov_inst_mult_238_n75, sec_nov_inst_mult_238_n74, 
      sec_nov_inst_mult_238_n73, sec_nov_inst_mult_238_n72, 
      sec_nov_inst_mult_238_n71, sec_nov_inst_mult_238_n70, 
      sec_nov_inst_mult_238_n69, sec_nov_inst_mult_238_n68, 
      sec_nov_inst_mult_238_n67, sec_nov_inst_mult_238_n65, 
      sec_nov_inst_mult_238_n64, sec_nov_inst_mult_238_n63, 
      sec_nov_inst_mult_238_n62, sec_nov_inst_mult_238_n60, 
      sec_nov_inst_mult_238_n59, sec_nov_inst_mult_238_n58, 
      sec_nov_inst_mult_238_n57, sec_nov_inst_mult_238_n56, 
      sec_nov_inst_mult_238_n55, sec_nov_inst_mult_238_n54, 
      sec_nov_inst_mult_238_n53, sec_nov_inst_mult_238_n52, 
      sec_nov_inst_mult_238_n51, sec_nov_inst_mult_238_n50, 
      sec_nov_inst_mult_238_n49, sec_nov_inst_mult_238_n48, 
      sec_nov_inst_mult_238_n47, sec_nov_inst_mult_238_n46, 
      sec_nov_inst_mult_238_n45, sec_nov_inst_mult_238_n44, 
      sec_nov_inst_mult_238_n43, sec_nov_inst_mult_238_n42, 
      sec_nov_inst_mult_238_n41, sec_nov_inst_mult_238_n40, 
      sec_nov_inst_mult_238_n39, sec_nov_inst_mult_238_n38, 
      sec_nov_inst_mult_238_n37, sec_nov_inst_mult_238_n36, 
      sec_nov_inst_mult_238_n35, sec_nov_inst_mult_238_n34, 
      sec_nov_inst_mult_238_n33, sec_nov_inst_mult_238_n31, 
      sec_nov_inst_mult_238_n30, sec_nov_inst_mult_238_n29, 
      sec_nov_inst_mult_238_n28, sec_nov_inst_mult_238_n27, 
      sec_nov_inst_mult_238_n26, sec_nov_inst_mult_238_n25, 
      sec_nov_inst_mult_238_n24, sec_nov_inst_mult_238_n23, 
      sec_nov_inst_mult_238_n21, sec_nov_inst_mult_238_n20, 
      sec_nov_inst_mult_238_n19, sec_nov_inst_mult_238_n18, 
      sec_nov_inst_mult_238_n17, sec_nov_inst_mult_238_n16, 
      sec_nov_inst_mult_238_n14, sec_nov_inst_mult_238_n13, 
      sec_nov_inst_mult_238_n12, sec_nov_inst_mult_238_n11, 
      sec_nov_inst_mult_238_n10, sec_nov_inst_mult_238_n9, 
      sec_nov_inst_mult_238_n8, sec_nov_inst_mult_238_n7, 
      sec_nov_inst_mult_238_n6, sec_nov_inst_mult_238_n5, 
      sec_nov_inst_mult_238_n4, sec_nov_inst_mult_238_n3, 
      sec_nov_inst_mult_238_n2 : std_logic;

begin
   
   sec_nov_inst_U152 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_arx_r1_reg_7_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, B => 
                           sec_nov_inst_n17, Z => sec_nov_inst_m_in_r_7_port);
   sec_nov_inst_U151 : AOI22D1 port map( A1 => sec_nov_inst_arx_d2_reg_7_port, 
                           A2 => sec_nov_inst_n16, B1 => 
                           sec_nov_inst_arx_d1_reg_7_port, B2 => 
                           sec_nov_inst_n15, Z => sec_nov_inst_n17);
   sec_nov_inst_U150 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_arx_r1_reg_6_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, B => 
                           sec_nov_inst_n14, Z => sec_nov_inst_m_in_r_6_port);
   sec_nov_inst_U149 : AOI22D1 port map( A1 => sec_nov_inst_arx_d2_reg_6_port, 
                           A2 => sec_nov_inst_n16, B1 => 
                           sec_nov_inst_arx_d1_reg_6_port, B2 => 
                           sec_nov_inst_n15, Z => sec_nov_inst_n14);
   sec_nov_inst_U148 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_arx_r1_reg_5_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, B => 
                           sec_nov_inst_n13, Z => sec_nov_inst_m_in_r_5_port);
   sec_nov_inst_U147 : AOI22D1 port map( A1 => sec_nov_inst_arx_d2_reg_5_port, 
                           A2 => sec_nov_inst_n16, B1 => 
                           sec_nov_inst_arx_d1_reg_5_port, B2 => 
                           sec_nov_inst_n15, Z => sec_nov_inst_n13);
   sec_nov_inst_U146 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_arx_r1_reg_4_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, B => 
                           sec_nov_inst_n12, Z => sec_nov_inst_m_in_r_4_port);
   sec_nov_inst_U145 : AOI22D1 port map( A1 => sec_nov_inst_arx_d2_reg_4_port, 
                           A2 => sec_nov_inst_n16, B1 => 
                           sec_nov_inst_arx_d1_reg_4_port, B2 => 
                           sec_nov_inst_n15, Z => sec_nov_inst_n12);
   sec_nov_inst_U144 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_arx_r1_reg_3_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, B => 
                           sec_nov_inst_n11, Z => sec_nov_inst_m_in_r_3_port);
   sec_nov_inst_U143 : AOI22D1 port map( A1 => sec_nov_inst_arx_d2_reg_3_port, 
                           A2 => sec_nov_inst_n16, B1 => 
                           sec_nov_inst_arx_d1_reg_3_port, B2 => 
                           sec_nov_inst_n15, Z => sec_nov_inst_n11);
   sec_nov_inst_U142 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_arx_r1_reg_2_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, B => 
                           sec_nov_inst_n10, Z => sec_nov_inst_m_in_r_2_port);
   sec_nov_inst_U141 : AOI22D1 port map( A1 => sec_nov_inst_arx_d2_reg_2_port, 
                           A2 => sec_nov_inst_n16, B1 => 
                           sec_nov_inst_arx_d1_reg_2_port, B2 => 
                           sec_nov_inst_n15, Z => sec_nov_inst_n10);
   sec_nov_inst_U140 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_arx_r1_reg_1_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, B => 
                           sec_nov_inst_n9, Z => sec_nov_inst_m_in_r_1_port);
   sec_nov_inst_U139 : AOI22D1 port map( A1 => sec_nov_inst_arx_d2_reg_1_port, 
                           A2 => sec_nov_inst_n16, B1 => 
                           sec_nov_inst_arx_d1_reg_1_port, B2 => 
                           sec_nov_inst_n15, Z => sec_nov_inst_n9);
   sec_nov_inst_U138 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_arx_r1_reg_0_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, B => 
                           sec_nov_inst_n8, Z => sec_nov_inst_m_in_r_0_port);
   sec_nov_inst_U137 : AOI22D1 port map( A1 => sec_nov_inst_arx_d2_reg_0_port, 
                           A2 => sec_nov_inst_n16, B1 => 
                           sec_nov_inst_arx_d1_reg_0_port, B2 => 
                           sec_nov_inst_n15, Z => sec_nov_inst_n8);
   sec_nov_inst_U136 : NOR2M1D1 port map( A1 => 
                           sec_nov_inst_arx_state_reg_1_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, Z => 
                           sec_nov_inst_n15);
   sec_nov_inst_U135 : NOR2D1 port map( A1 => sec_nov_inst_arx_state_reg_3_port
                           , A2 => sec_nov_inst_arx_state_reg_1_port, Z => 
                           sec_nov_inst_n16);
   sec_nov_inst_U134 : EXOR2D1 port map( A1 => sec_nov_inst_N123, A2 => 
                           sec_nov_inst_N124, Z => sec_nov_inst_a_out_0_port);
   sec_nov_inst_U133 : AND2D1 port map( A1 => sec_nov_inst_N124, A2 => 
                           sec_nov_inst_N123, Z => 
                           sec_nov_inst_add_416_C239_rn_carry_1_port);
   sec_nov_inst_U132 : EXOR2D1 port map( A1 => sec_nov_inst_N125, A2 => 
                           sec_nov_inst_add_416_C239_rn_carry_1_port, Z => 
                           sec_nov_inst_a_out_1_port);
   sec_nov_inst_U131 : AND2D1 port map( A1 => 
                           sec_nov_inst_add_416_C239_rn_carry_1_port, A2 => 
                           sec_nov_inst_N125, Z => 
                           sec_nov_inst_add_416_C239_rn_carry_2_port);
   sec_nov_inst_U130 : EXOR2D1 port map( A1 => sec_nov_inst_N126, A2 => 
                           sec_nov_inst_add_416_C239_rn_carry_2_port, Z => 
                           sec_nov_inst_a_out_2_port);
   sec_nov_inst_U129 : AND2D1 port map( A1 => 
                           sec_nov_inst_add_416_C239_rn_carry_2_port, A2 => 
                           sec_nov_inst_N126, Z => 
                           sec_nov_inst_add_416_C239_rn_carry_3_port);
   sec_nov_inst_U128 : EXOR2D1 port map( A1 => sec_nov_inst_N127, A2 => 
                           sec_nov_inst_add_416_C239_rn_carry_3_port, Z => 
                           sec_nov_inst_a_out_3_port);
   sec_nov_inst_U127 : AND2D1 port map( A1 => 
                           sec_nov_inst_add_416_C239_rn_carry_3_port, A2 => 
                           sec_nov_inst_N127, Z => 
                           sec_nov_inst_add_416_C239_rn_carry_4_port);
   sec_nov_inst_U126 : EXOR2D1 port map( A1 => sec_nov_inst_N128, A2 => 
                           sec_nov_inst_add_416_C239_rn_carry_4_port, Z => 
                           sec_nov_inst_a_out_4_port);
   sec_nov_inst_U125 : AND2D1 port map( A1 => 
                           sec_nov_inst_add_416_C239_rn_carry_4_port, A2 => 
                           sec_nov_inst_N128, Z => 
                           sec_nov_inst_add_416_C239_rn_carry_5_port);
   sec_nov_inst_U124 : EXOR2D1 port map( A1 => sec_nov_inst_N129, A2 => 
                           sec_nov_inst_add_416_C239_rn_carry_5_port, Z => 
                           sec_nov_inst_a_out_5_port);
   sec_nov_inst_U123 : AND2D1 port map( A1 => 
                           sec_nov_inst_add_416_C239_rn_carry_5_port, A2 => 
                           sec_nov_inst_N129, Z => 
                           sec_nov_inst_add_416_C239_rn_carry_6_port);
   sec_nov_inst_U122 : EXOR2D1 port map( A1 => sec_nov_inst_N130, A2 => 
                           sec_nov_inst_add_416_C239_rn_carry_6_port, Z => 
                           sec_nov_inst_a_out_6_port);
   sec_nov_inst_U121 : AND2D1 port map( A1 => 
                           sec_nov_inst_add_416_C239_rn_carry_6_port, A2 => 
                           sec_nov_inst_N130, Z => 
                           sec_nov_inst_add_416_C239_rn_carry_7_port);
   sec_nov_inst_U120 : EXOR2D1 port map( A1 => sec_nov_inst_N131, A2 => 
                           sec_nov_inst_add_416_C239_rn_carry_7_port, Z => 
                           sec_nov_inst_a_out_7_port);
   sec_nov_inst_U119 : TIELO port map( Z => sec_nov_inst_n7);
   sec_nov_inst_U118 : INVD1 port map( A => resetn, Z => sec_nov_inst_n6);
   sec_nov_inst_U117 : INVD1 port map( A => sec_nov_inst_n6, Z => 
                           sec_nov_inst_n2);
   sec_nov_inst_U98 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_14_port, Z 
                           => sec_nov_inst_n39);
   sec_nov_inst_U97 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_13_port, Z 
                           => sec_nov_inst_n25);
   sec_nov_inst_U96 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_12_port, Z 
                           => sec_nov_inst_n26);
   sec_nov_inst_U95 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_11_port, Z 
                           => sec_nov_inst_n27);
   sec_nov_inst_U94 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_10_port, Z 
                           => sec_nov_inst_n28);
   sec_nov_inst_U93 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_9_port, Z =>
                           sec_nov_inst_n29);
   sec_nov_inst_U92 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_8_port, Z =>
                           sec_nov_inst_n30);
   sec_nov_inst_U91 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_14_port, Z 
                           => sec_nov_inst_n24);
   sec_nov_inst_U90 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_7_port, Z =>
                           sec_nov_inst_n31);
   sec_nov_inst_U89 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_6_port, Z =>
                           sec_nov_inst_n32);
   sec_nov_inst_U88 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_6_port, Z =>
                           sec_nov_inst_n47);
   sec_nov_inst_U87 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_4_port, Z =>
                           sec_nov_inst_n49);
   sec_nov_inst_U86 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_4_port, Z =>
                           sec_nov_inst_n34);
   sec_nov_inst_U85 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_3_port, Z =>
                           sec_nov_inst_n50);
   sec_nov_inst_U84 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_3_port, Z =>
                           sec_nov_inst_n35);
   sec_nov_inst_U83 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_2_port, Z =>
                           sec_nov_inst_n51);
   sec_nov_inst_U82 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_2_port, Z =>
                           sec_nov_inst_n36);
   sec_nov_inst_U81 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_0_port, Z =>
                           sec_nov_inst_n85);
   sec_nov_inst_U80 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_1_port, Z =>
                           sec_nov_inst_n58);
   sec_nov_inst_U79 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_5_port, Z =>
                           sec_nov_inst_n33);
   sec_nov_inst_U78 : NOR2D1 port map( A1 => sec_nov_inst_n78, A2 => 
                           sec_nov_inst_n33, Z => sec_nov_inst_a_in_l_5_port);
   sec_nov_inst_U77 : NAN3D1 port map( A1 => sec_nov_inst_arx_state_reg_1_port,
                           A2 => sec_nov_inst_arx_state_reg_0_port, A3 => 
                           sec_nov_inst_n84, Z => sec_nov_inst_n54);
   sec_nov_inst_U76 : NOR2D1 port map( A1 => sec_nov_inst_arx_state_reg_0_port,
                           A2 => sec_nov_inst_arx_state_reg_1_port, Z => 
                           sec_nov_inst_n83);
   sec_nov_inst_U75 : NAN3D1 port map( A1 => sec_nov_inst_arx_state_reg_0_port,
                           A2 => sec_nov_inst_n80, A3 => 
                           sec_nov_inst_arx_state_reg_1_port, Z => 
                           sec_nov_inst_n53);
   sec_nov_inst_U74 : NOR2M1D1 port map( A1 => 
                           sec_nov_inst_arx_state_reg_2_port, A2 => 
                           sec_nov_inst_arx_state_reg_3_port, Z => 
                           sec_nov_inst_n80);
   sec_nov_inst_U73 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_0_port, Z =>
                           sec_nov_inst_n38);
   sec_nov_inst_U72 : NOR2D1 port map( A1 => sec_nov_inst_n78, A2 => 
                           sec_nov_inst_n38, Z => sec_nov_inst_a_in_l_0_port);
   sec_nov_inst_U71 : NOR2D1 port map( A1 => sec_nov_inst_arx_state_reg_2_port,
                           A2 => sec_nov_inst_arx_state_reg_3_port, Z => 
                           sec_nov_inst_n84);
   sec_nov_inst_U70 : NOR2M1D1 port map( A1 => 
                           sec_nov_inst_arx_state_reg_1_port, A2 => 
                           sec_nov_inst_arx_state_reg_0_port, Z => 
                           sec_nov_inst_n81);
   sec_nov_inst_U69 : INVD1 port map( A => sec_nov_inst_arx_r2_reg_1_port, Z =>
                           sec_nov_inst_n37);
   sec_nov_inst_U68 : NOR2D1 port map( A1 => sec_nov_inst_n78, A2 => 
                           sec_nov_inst_n37, Z => sec_nov_inst_a_in_l_1_port);
   sec_nov_inst_U67 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_13_port, Z 
                           => sec_nov_inst_n40);
   sec_nov_inst_U66 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_12_port, Z 
                           => sec_nov_inst_n41);
   sec_nov_inst_U65 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_11_port, Z 
                           => sec_nov_inst_n42);
   sec_nov_inst_U64 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_10_port, Z 
                           => sec_nov_inst_n43);
   sec_nov_inst_U63 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_9_port, Z =>
                           sec_nov_inst_n44);
   sec_nov_inst_U62 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_8_port, Z =>
                           sec_nov_inst_n45);
   sec_nov_inst_U61 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_7_port, Z =>
                           sec_nov_inst_n46);
   sec_nov_inst_U60 : INVD1 port map( A => sec_nov_inst_arx_r3_reg_5_port, Z =>
                           sec_nov_inst_n48);
   sec_nov_inst_U59 : NOR2D1 port map( A1 => sec_nov_inst_n76, A2 => 
                           sec_nov_inst_n48, Z => sec_nov_inst_a_in_r_5_port);
   sec_nov_inst_U58 : NOR2M1D1 port map( A1 => 
                           sec_nov_inst_arx_state_reg_0_port, A2 => 
                           sec_nov_inst_arx_state_reg_1_port, Z => 
                           sec_nov_inst_n79);
   sec_nov_inst_U57 : NOR2M1D1 port map( A1 => 
                           sec_nov_inst_arx_state_reg_3_port, A2 => 
                           sec_nov_inst_arx_state_reg_2_port, Z => 
                           sec_nov_inst_n82);
   sec_nov_inst_U56 : INVD1 port map( A => sec_nov_inst_n6, Z => 
                           sec_nov_inst_n5);
   sec_nov_inst_U55 : INVD1 port map( A => sec_nov_inst_n6, Z => 
                           sec_nov_inst_n4);
   sec_nov_inst_U54 : INVD1 port map( A => sec_nov_inst_n6, Z => 
                           sec_nov_inst_n3);
   sec_nov_inst_U53 : NAN4D1 port map( A1 => sec_nov_inst_n54, A2 => 
                           sec_nov_inst_n55, A3 => sec_nov_inst_n56, A4 => 
                           sec_nov_inst_n57, Z => sec_nov_inst_state_2_port);
   sec_nov_inst_U52 : NAN2D1 port map( A1 => sec_nov_inst_n52, A2 => 
                           sec_nov_inst_n53, Z => sec_nov_inst_state_3_port);
   sec_nov_inst_U51 : AND3D1 port map( A1 => sec_nov_inst_n54, A2 => 
                           sec_nov_inst_n53, A3 => sec_nov_inst_n67, Z => 
                           sec_nov_inst_n65);
   sec_nov_inst_U50 : NAN2D1 port map( A1 => sec_nov_inst_n84, A2 => 
                           sec_nov_inst_n81, Z => sec_nov_inst_n69);
   sec_nov_inst_U49 : NAN2D1 port map( A1 => sec_nov_inst_n83, A2 => 
                           sec_nov_inst_n80, Z => sec_nov_inst_n55);
   sec_nov_inst_U48 : NAN2D1 port map( A1 => sec_nov_inst_n79, A2 => 
                           sec_nov_inst_n80, Z => sec_nov_inst_n56);
   sec_nov_inst_U47 : NAN2D1 port map( A1 => sec_nov_inst_n84, A2 => 
                           sec_nov_inst_n83, Z => sec_nov_inst_n64);
   sec_nov_inst_U46 : NAN2D1 port map( A1 => sec_nov_inst_n81, A2 => 
                           sec_nov_inst_n82, Z => sec_nov_inst_n67);
   sec_nov_inst_U45 : AND2D1 port map( A1 => sec_nov_inst_n53, A2 => 
                           sec_nov_inst_n57, Z => sec_nov_inst_n74);
   sec_nov_inst_U44 : NAN2D1 port map( A1 => sec_nov_inst_n81, A2 => 
                           sec_nov_inst_n80, Z => sec_nov_inst_n57);
   sec_nov_inst_U43 : NOR2D1 port map( A1 => sec_nov_inst_n78, A2 => 
                           sec_nov_inst_n34, Z => sec_nov_inst_a_in_l_4_port);
   sec_nov_inst_U42 : NOR2D1 port map( A1 => sec_nov_inst_n76, A2 => 
                           sec_nov_inst_n49, Z => sec_nov_inst_a_in_r_4_port);
   sec_nov_inst_U41 : NOR2D1 port map( A1 => sec_nov_inst_n78, A2 => 
                           sec_nov_inst_n35, Z => sec_nov_inst_a_in_l_3_port);
   sec_nov_inst_U40 : NOR2D1 port map( A1 => sec_nov_inst_n76, A2 => 
                           sec_nov_inst_n50, Z => sec_nov_inst_a_in_r_3_port);
   sec_nov_inst_U39 : NOR2D1 port map( A1 => sec_nov_inst_n78, A2 => 
                           sec_nov_inst_n36, Z => sec_nov_inst_a_in_l_2_port);
   sec_nov_inst_U38 : NOR2D1 port map( A1 => sec_nov_inst_n76, A2 => 
                           sec_nov_inst_n51, Z => sec_nov_inst_a_in_r_2_port);
   sec_nov_inst_U37 : NOR2D1 port map( A1 => sec_nov_inst_n78, A2 => 
                           sec_nov_inst_n32, Z => sec_nov_inst_a_in_l_6_port);
   sec_nov_inst_U36 : NOR2D1 port map( A1 => sec_nov_inst_n76, A2 => 
                           sec_nov_inst_n47, Z => sec_nov_inst_a_in_r_6_port);
   sec_nov_inst_U35 : NAN2D1 port map( A1 => sec_nov_inst_n84, A2 => 
                           sec_nov_inst_n79, Z => sec_nov_inst_n62);
   sec_nov_inst_U34 : NAN3D1 port map( A1 => sec_nov_inst_n54, A2 => 
                           sec_nov_inst_n22, A3 => sec_nov_inst_n69, Z => 
                           sec_nov_inst_m_in_l_6_port);
   sec_nov_inst_U33 : NOR2D1 port map( A1 => sec_nov_inst_n76, A2 => 
                           sec_nov_inst_n58, Z => sec_nov_inst_a_in_r_1_port);
   sec_nov_inst_U32 : NOR2D1 port map( A1 => sec_nov_inst_n76, A2 => 
                           sec_nov_inst_n85, Z => sec_nov_inst_a_in_r_0_port);
   sec_nov_inst_U31 : NAN2D1 port map( A1 => sec_nov_inst_n83, A2 => 
                           sec_nov_inst_n82, Z => sec_nov_inst_n71);
   sec_nov_inst_U30 : NAN2D1 port map( A1 => sec_nov_inst_n79, A2 => 
                           sec_nov_inst_n82, Z => sec_nov_inst_n63);
   sec_nov_inst_U29 : NAN3D1 port map( A1 => sec_nov_inst_n64, A2 => 
                           sec_nov_inst_n23, A3 => sec_nov_inst_n65, Z => 
                           sec_nov_inst_n61);
   sec_nov_inst_U28 : AND3D1 port map( A1 => sec_nov_inst_n56, A2 => 
                           sec_nov_inst_n63, A3 => sec_nov_inst_n57, Z => 
                           sec_nov_inst_n73);
   sec_nov_inst_U27 : NAN3D1 port map( A1 => sec_nov_inst_n62, A2 => 
                           sec_nov_inst_n69, A3 => sec_nov_inst_n73, Z => 
                           sec_nov_inst_state_1_port);
   sec_nov_inst_U26 : NAN4D1 port map( A1 => sec_nov_inst_n65, A2 => 
                           sec_nov_inst_n55, A3 => sec_nov_inst_n71, A4 => 
                           sec_nov_inst_n23, Z => sec_nov_inst_n72);
   sec_nov_inst_U25 : NAN3D1 port map( A1 => sec_nov_inst_n67, A2 => 
                           sec_nov_inst_n56, A3 => sec_nov_inst_n59, Z => 
                           sec_nov_inst_n66);
   sec_nov_inst_U24 : NAN2D1 port map( A1 => sec_nov_inst_n65, A2 => 
                           sec_nov_inst_n20, Z => sec_nov_inst_n68);
   sec_nov_inst_U23 : INVD1 port map( A => sec_nov_inst_n68, Z => 
                           sec_nov_inst_n19);
   sec_nov_inst_U22 : NAN3D1 port map( A1 => sec_nov_inst_n62, A2 => 
                           sec_nov_inst_n63, A3 => sec_nov_inst_n19, Z => 
                           sec_nov_inst_n60);
   sec_nov_inst_U21 : AND3D1 port map( A1 => sec_nov_inst_n63, A2 => 
                           sec_nov_inst_n20, A3 => sec_nov_inst_n62, Z => 
                           sec_nov_inst_n59);
   sec_nov_inst_U20 : AND3D1 port map( A1 => sec_nov_inst_n57, A2 => 
                           sec_nov_inst_n64, A3 => sec_nov_inst_n71, Z => 
                           sec_nov_inst_n70);
   sec_nov_inst_U19 : NAN3D1 port map( A1 => sec_nov_inst_n69, A2 => 
                           sec_nov_inst_n55, A3 => sec_nov_inst_n70, Z => 
                           sec_nov_inst_state_0_port);
   sec_nov_inst_U18 : AND2D1 port map( A1 => sec_nov_inst_n77, A2 => 
                           sec_nov_inst_n67, Z => sec_nov_inst_n75);
   sec_nov_inst_U17 : AND2D1 port map( A1 => sec_nov_inst_n74, A2 => 
                           sec_nov_inst_n56, Z => sec_nov_inst_n77);
   sec_nov_inst_U16 : NAN2D1 port map( A1 => sec_nov_inst_n74, A2 => 
                           sec_nov_inst_n22, Z => sec_nov_inst_m_in_l_7_port);
   sec_nov_inst_U15 : INVD1 port map( A => sec_nov_inst_m_in_l_6_port, Z => 
                           sec_nov_inst_n21);
   sec_nov_inst_U14 : NAN2D1 port map( A1 => sec_nov_inst_n64, A2 => 
                           sec_nov_inst_n62, Z => sec_nov_inst_m_in_l_2_port);
   sec_nov_inst_U13 : AND2D1 port map( A1 => sec_nov_inst_n76, A2 => 
                           sec_nov_inst_n67, Z => sec_nov_inst_n78);
   sec_nov_inst_U12 : AND3D1 port map( A1 => sec_nov_inst_n55, A2 => 
                           sec_nov_inst_n21, A3 => sec_nov_inst_n52, Z => 
                           sec_nov_inst_n76);
   sec_nov_inst_U11 : NAN2D1 port map( A1 => sec_nov_inst_n74, A2 => 
                           sec_nov_inst_n18, Z => sec_nov_inst_m_in_l_4_port);
   sec_nov_inst_U10 : AND2D1 port map( A1 => sec_nov_inst_n63, A2 => 
                           sec_nov_inst_n71, Z => sec_nov_inst_n52);
   sec_nov_inst_U9 : NAN4D1 port map( A1 => sec_nov_inst_n52, A2 => 
                           sec_nov_inst_n67, A3 => sec_nov_inst_n55, A4 => 
                           sec_nov_inst_n56, Z => sec_nov_inst_m_in_l_5_port);
   sec_nov_inst_U8 : INVD1 port map( A => sec_nov_inst_state_1_port, Z => 
                           sec_nov_inst_n23);
   sec_nov_inst_U7 : INVD1 port map( A => sec_nov_inst_state_0_port, Z => 
                           sec_nov_inst_n20);
   sec_nov_inst_U6 : NAN2D1 port map( A1 => sec_nov_inst_n18, A2 => 
                           sec_nov_inst_n21, Z => sec_nov_inst_m_in_l_0_port);
   sec_nov_inst_U5 : INVD1 port map( A => sec_nov_inst_m_in_l_2_port, Z => 
                           sec_nov_inst_n22);
   sec_nov_inst_U4 : INVD1 port map( A => sec_nov_inst_m_in_l_5_port, Z => 
                           sec_nov_inst_n18);
   sec_nov_inst_U3 : NAN4D1 port map( A1 => sec_nov_inst_n59, A2 => 
                           sec_nov_inst_n54, A3 => sec_nov_inst_n56, A4 => 
                           sec_nov_inst_n53, Z => sec_nov_inst_n1);
   sec_nov_inst_arx_d0_reg_reg_0 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_0_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n3, Q => 
                           sec_nov_inst_arx_d0_reg_0_port);
   sec_nov_inst_arx_d0_reg_reg_1 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_1_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n3, Q => 
                           sec_nov_inst_arx_d0_reg_1_port);
   sec_nov_inst_arx_d0_reg_reg_2 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_2_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_d0_reg_2_port);
   sec_nov_inst_arx_d0_reg_reg_3 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_3_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_d0_reg_3_port);
   sec_nov_inst_arx_d0_reg_reg_4 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_4_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_d0_reg_4_port);
   sec_nov_inst_arx_d0_reg_reg_5 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_5_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_d0_reg_5_port);
   sec_nov_inst_arx_d0_reg_reg_6 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_6_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_d0_reg_6_port);
   sec_nov_inst_arx_o1_reg_reg_0 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_0_port, CEB => sec_nov_inst_n1, 
                           CK => clock, RB => sec_nov_inst_n2, Q => data_out(0)
                           );
   sec_nov_inst_arx_o1_reg_reg_1 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_1_port, CEB => sec_nov_inst_n1, 
                           CK => clock, RB => sec_nov_inst_n2, Q => data_out(1)
                           );
   sec_nov_inst_arx_o1_reg_reg_2 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_2_port, CEB => sec_nov_inst_n1, 
                           CK => clock, RB => sec_nov_inst_n2, Q => data_out(2)
                           );
   sec_nov_inst_arx_o1_reg_reg_3 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_3_port, CEB => sec_nov_inst_n1, 
                           CK => clock, RB => sec_nov_inst_n2, Q => data_out(3)
                           );
   sec_nov_inst_arx_o1_reg_reg_4 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_4_port, CEB => sec_nov_inst_n1, 
                           CK => clock, RB => sec_nov_inst_n2, Q => data_out(4)
                           );
   sec_nov_inst_arx_o1_reg_reg_5 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_5_port, CEB => sec_nov_inst_n1, 
                           CK => clock, RB => sec_nov_inst_n2, Q => data_out(5)
                           );
   sec_nov_inst_arx_o1_reg_reg_6 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_6_port, CEB => sec_nov_inst_n1, 
                           CK => clock, RB => sec_nov_inst_n2, Q => data_out(6)
                           );
   sec_nov_inst_arx_o1_reg_reg_7 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_7_port, CEB => sec_nov_inst_n1, 
                           CK => clock, RB => sec_nov_inst_n2, Q => data_out(7)
                           );
   sec_nov_inst_arx_d0_reg_reg_7 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_7_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_d0_reg_7_port);
   sec_nov_inst_arx_state_reg_reg_3 : DFFRPQ1 port map( D => 
                           sec_nov_inst_state_3_port, CK => clock, RB => resetn
                           , Q => sec_nov_inst_arx_state_reg_3_port);
   sec_nov_inst_arx_state_reg_reg_0 : DFFRPQ1 port map( D => 
                           sec_nov_inst_state_0_port, CK => clock, RB => resetn
                           , Q => sec_nov_inst_arx_state_reg_0_port);
   sec_nov_inst_arx_state_reg_reg_1 : DFFRPQ1 port map( D => 
                           sec_nov_inst_state_1_port, CK => clock, RB => resetn
                           , Q => sec_nov_inst_arx_state_reg_1_port);
   sec_nov_inst_arx_state_reg_reg_2 : DFFRPQ1 port map( D => 
                           sec_nov_inst_state_2_port, CK => clock, RB => resetn
                           , Q => sec_nov_inst_arx_state_reg_2_port);
   sec_nov_inst_arx_d2_reg_reg_1 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d1_reg_1_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n2,
                           Q => sec_nov_inst_arx_d2_reg_1_port);
   sec_nov_inst_arx_d1_reg_reg_1 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d0_reg_1_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d1_reg_1_port);
   sec_nov_inst_arx_d2_reg_reg_0 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d1_reg_0_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n2,
                           Q => sec_nov_inst_arx_d2_reg_0_port);
   sec_nov_inst_arx_d1_reg_reg_0 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d0_reg_0_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d1_reg_0_port);
   sec_nov_inst_arx_r1_reg_reg_0 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_0_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r1_reg_0_port);
   sec_nov_inst_arx_r1_reg_reg_1 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_1_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r1_reg_1_port);
   sec_nov_inst_arx_d2_reg_reg_3 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d1_reg_3_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n2,
                           Q => sec_nov_inst_arx_d2_reg_3_port);
   sec_nov_inst_arx_d1_reg_reg_3 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d0_reg_3_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d1_reg_3_port);
   sec_nov_inst_arx_d2_reg_reg_2 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d1_reg_2_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n2,
                           Q => sec_nov_inst_arx_d2_reg_2_port);
   sec_nov_inst_arx_r1_reg_reg_3 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_3_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r1_reg_3_port);
   sec_nov_inst_arx_d1_reg_reg_2 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d0_reg_2_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d1_reg_2_port);
   sec_nov_inst_arx_r1_reg_reg_2 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_2_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r1_reg_2_port);
   sec_nov_inst_arx_d2_reg_reg_4 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d1_reg_4_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n2,
                           Q => sec_nov_inst_arx_d2_reg_4_port);
   sec_nov_inst_arx_d1_reg_reg_4 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d0_reg_4_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d1_reg_4_port);
   sec_nov_inst_arx_r1_reg_reg_4 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_4_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r1_reg_4_port);
   sec_nov_inst_arx_d2_reg_reg_5 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d1_reg_5_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d2_reg_5_port);
   sec_nov_inst_arx_d1_reg_reg_5 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d0_reg_5_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d1_reg_5_port);
   sec_nov_inst_arx_r1_reg_reg_5 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_5_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_r1_reg_5_port);
   sec_nov_inst_arx_r3_reg_reg_1 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_1_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r3_reg_1_port);
   sec_nov_inst_arx_r2_reg_reg_1 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_1_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_1_port);
   sec_nov_inst_arx_d2_reg_reg_6 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d1_reg_6_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d2_reg_6_port);
   sec_nov_inst_arx_d1_reg_reg_6 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d0_reg_6_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d1_reg_6_port);
   sec_nov_inst_arx_r2_reg_reg_0 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_0_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_0_port);
   sec_nov_inst_arx_r1_reg_reg_6 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_6_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_r1_reg_6_port);
   sec_nov_inst_arx_r3_reg_reg_0 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_0_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r3_reg_0_port);
   sec_nov_inst_arx_r2_reg_reg_2 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_2_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_2_port);
   sec_nov_inst_arx_r3_reg_reg_2 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_2_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r3_reg_2_port);
   sec_nov_inst_arx_d2_reg_reg_7 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d1_reg_7_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d2_reg_7_port);
   sec_nov_inst_arx_d1_reg_reg_7 : DFERPQ1 port map( D => 
                           sec_nov_inst_arx_d0_reg_7_port, CEB => 
                           sec_nov_inst_n1, CK => clock, RB => sec_nov_inst_n3,
                           Q => sec_nov_inst_arx_d1_reg_7_port);
   sec_nov_inst_arx_r1_reg_reg_7 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_7_port, CEB => sec_nov_inst_n60, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_r1_reg_7_port);
   sec_nov_inst_arx_r2_reg_reg_3 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_3_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_3_port);
   sec_nov_inst_arx_r3_reg_reg_3 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_3_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r3_reg_3_port);
   sec_nov_inst_arx_r2_reg_reg_4 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_4_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_4_port);
   sec_nov_inst_arx_r3_reg_reg_4 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_4_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_4_port);
   sec_nov_inst_arx_r2_reg_reg_5 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_5_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_5_port);
   sec_nov_inst_arx_r3_reg_reg_5 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_5_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_5_port);
   sec_nov_inst_arx_r3_reg_reg_6 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_6_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_6_port);
   sec_nov_inst_arx_r2_reg_reg_6 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_6_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_6_port);
   sec_nov_inst_arx_r4_reg_reg_0 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_0_port, CEB => sec_nov_inst_n61, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r4_reg_0_port);
   sec_nov_inst_arx_i1_reg_reg_0 : DFERPQ1 port map( D => data_in(0), CEB => 
                           sec_nov_inst_n72, CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_i1_reg_0_port);
   sec_nov_inst_arx_r3_reg_reg_7 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_7_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_7_port);
   sec_nov_inst_arx_r2_reg_reg_7 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_7_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_7_port);
   sec_nov_inst_arx_r4_reg_reg_1 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_1_port, CEB => sec_nov_inst_n61, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r4_reg_1_port);
   sec_nov_inst_arx_i1_reg_reg_1 : DFERPQ1 port map( D => data_in(1), CEB => 
                           sec_nov_inst_n72, CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_i1_reg_1_port);
   sec_nov_inst_arx_r3_reg_reg_8 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_8_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_8_port);
   sec_nov_inst_arx_r2_reg_reg_8 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_8_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_8_port);
   sec_nov_inst_arx_r4_reg_reg_2 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_2_port, CEB => sec_nov_inst_n61, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r4_reg_2_port);
   sec_nov_inst_arx_i1_reg_reg_2 : DFERPQ1 port map( D => data_in(2), CEB => 
                           sec_nov_inst_n72, CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_i1_reg_2_port);
   sec_nov_inst_arx_r3_reg_reg_9 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_9_port, CEB => sec_nov_inst_n66, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_9_port);
   sec_nov_inst_arx_r2_reg_reg_9 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_9_port, CEB => sec_nov_inst_n68, 
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_9_port);
   sec_nov_inst_arx_r4_reg_reg_3 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_3_port, CEB => sec_nov_inst_n61, 
                           CK => clock, RB => sec_nov_inst_n5, Q => 
                           sec_nov_inst_arx_r4_reg_3_port);
   sec_nov_inst_arx_i1_reg_reg_3 : DFERPQ1 port map( D => data_in(3), CEB => 
                           sec_nov_inst_n72, CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_i1_reg_3_port);
   sec_nov_inst_arx_r3_reg_reg_10 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_10_port, CEB => sec_nov_inst_n66,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_10_port);
   sec_nov_inst_arx_r2_reg_reg_10 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_10_port, CEB => sec_nov_inst_n68,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_10_port);
   sec_nov_inst_arx_r4_reg_reg_4 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_4_port, CEB => sec_nov_inst_n61, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_r4_reg_4_port);
   sec_nov_inst_arx_i1_reg_reg_4 : DFERPQ1 port map( D => data_in(4), CEB => 
                           sec_nov_inst_n72, CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_i1_reg_4_port);
   sec_nov_inst_arx_r3_reg_reg_11 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_11_port, CEB => sec_nov_inst_n66,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_11_port);
   sec_nov_inst_arx_r2_reg_reg_11 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_11_port, CEB => sec_nov_inst_n68,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_11_port);
   sec_nov_inst_arx_r4_reg_reg_5 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_5_port, CEB => sec_nov_inst_n61, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_r4_reg_5_port);
   sec_nov_inst_arx_i1_reg_reg_5 : DFERPQ1 port map( D => data_in(5), CEB => 
                           sec_nov_inst_n72, CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_i1_reg_5_port);
   sec_nov_inst_arx_r3_reg_reg_12 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_12_port, CEB => sec_nov_inst_n66,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_12_port);
   sec_nov_inst_arx_r2_reg_reg_12 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_12_port, CEB => sec_nov_inst_n68,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_12_port);
   sec_nov_inst_arx_r4_reg_reg_6 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_6_port, CEB => sec_nov_inst_n61, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_r4_reg_6_port);
   sec_nov_inst_arx_i1_reg_reg_6 : DFERPQ1 port map( D => data_in(6), CEB => 
                           sec_nov_inst_n72, CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_i1_reg_6_port);
   sec_nov_inst_arx_r3_reg_reg_13 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_13_port, CEB => sec_nov_inst_n66,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_13_port);
   sec_nov_inst_arx_r2_reg_reg_13 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_13_port, CEB => sec_nov_inst_n68,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_13_port);
   sec_nov_inst_arx_r4_reg_reg_7 : DFERPQ1 port map( D => 
                           sec_nov_inst_a_out_7_port, CEB => sec_nov_inst_n61, 
                           CK => clock, RB => sec_nov_inst_n4, Q => 
                           sec_nov_inst_arx_r4_reg_7_port);
   sec_nov_inst_arx_i1_reg_reg_7 : DFERPQ1 port map( D => data_in(7), CEB => 
                           sec_nov_inst_n72, CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_i1_reg_7_port);
   sec_nov_inst_arx_r3_reg_reg_14 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_14_port, CEB => sec_nov_inst_n66,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r3_reg_14_port);
   sec_nov_inst_arx_r2_reg_reg_14 : DFERPQ1 port map( D => 
                           sec_nov_inst_m_out_14_port, CEB => sec_nov_inst_n68,
                           CK => clock, RB => resetn, Q => 
                           sec_nov_inst_arx_r2_reg_14_port);
   sec_nov_inst_U116 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_i1_reg_3_port, A2 => 
                           sec_nov_inst_n77, B1 => sec_nov_inst_n78, B2 => 
                           sec_nov_inst_n28, Z => sec_nov_inst_a_in_l_10_port);
   sec_nov_inst_U115 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_i1_reg_4_port, A2 => 
                           sec_nov_inst_n77, B1 => sec_nov_inst_n78, B2 => 
                           sec_nov_inst_n27, Z => sec_nov_inst_a_in_l_11_port);
   sec_nov_inst_U114 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_i1_reg_5_port, A2 => 
                           sec_nov_inst_n77, B1 => sec_nov_inst_n78, B2 => 
                           sec_nov_inst_n26, Z => sec_nov_inst_a_in_l_12_port);
   sec_nov_inst_U113 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_i1_reg_6_port, A2 => 
                           sec_nov_inst_n77, B1 => sec_nov_inst_n78, B2 => 
                           sec_nov_inst_n25, Z => sec_nov_inst_a_in_l_13_port);
   sec_nov_inst_U112 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_i1_reg_7_port, A2 => 
                           sec_nov_inst_n77, B1 => sec_nov_inst_n78, B2 => 
                           sec_nov_inst_n24, Z => sec_nov_inst_a_in_l_14_port);
   sec_nov_inst_U111 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_i1_reg_0_port, A2 => 
                           sec_nov_inst_n77, B1 => sec_nov_inst_n78, B2 => 
                           sec_nov_inst_n31, Z => sec_nov_inst_a_in_l_7_port);
   sec_nov_inst_U110 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_i1_reg_1_port, A2 => 
                           sec_nov_inst_n77, B1 => sec_nov_inst_n78, B2 => 
                           sec_nov_inst_n30, Z => sec_nov_inst_a_in_l_8_port);
   sec_nov_inst_U109 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_i1_reg_2_port, A2 => 
                           sec_nov_inst_n77, B1 => sec_nov_inst_n78, B2 => 
                           sec_nov_inst_n29, Z => sec_nov_inst_a_in_l_9_port);
   sec_nov_inst_U108 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_r4_reg_3_port, A2 => 
                           sec_nov_inst_n75, B1 => sec_nov_inst_n76, B2 => 
                           sec_nov_inst_n43, Z => sec_nov_inst_a_in_r_10_port);
   sec_nov_inst_U107 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_r4_reg_4_port, A2 => 
                           sec_nov_inst_n75, B1 => sec_nov_inst_n76, B2 => 
                           sec_nov_inst_n42, Z => sec_nov_inst_a_in_r_11_port);
   sec_nov_inst_U106 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_r4_reg_5_port, A2 => 
                           sec_nov_inst_n75, B1 => sec_nov_inst_n76, B2 => 
                           sec_nov_inst_n41, Z => sec_nov_inst_a_in_r_12_port);
   sec_nov_inst_U105 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_r4_reg_6_port, A2 => 
                           sec_nov_inst_n75, B1 => sec_nov_inst_n76, B2 => 
                           sec_nov_inst_n40, Z => sec_nov_inst_a_in_r_13_port);
   sec_nov_inst_U104 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_r4_reg_7_port, A2 => 
                           sec_nov_inst_n75, B1 => sec_nov_inst_n76, B2 => 
                           sec_nov_inst_n39, Z => sec_nov_inst_a_in_r_14_port);
   sec_nov_inst_U103 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_r4_reg_0_port, A2 => 
                           sec_nov_inst_n75, B1 => sec_nov_inst_n76, B2 => 
                           sec_nov_inst_n46, Z => sec_nov_inst_a_in_r_7_port);
   sec_nov_inst_U102 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_r4_reg_1_port, A2 => 
                           sec_nov_inst_n75, B1 => sec_nov_inst_n76, B2 => 
                           sec_nov_inst_n45, Z => sec_nov_inst_a_in_r_8_port);
   sec_nov_inst_U101 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_arx_r4_reg_2_port, A2 => 
                           sec_nov_inst_n75, B1 => sec_nov_inst_n76, B2 => 
                           sec_nov_inst_n44, Z => sec_nov_inst_a_in_r_9_port);
   sec_nov_inst_U100 : NAN3M1D1 port map( A1 => sec_nov_inst_m_in_l_7_port, A2 
                           => sec_nov_inst_n54, A3 => sec_nov_inst_n69, Z => 
                           sec_nov_inst_m_in_l_1_port);
   sec_nov_inst_U99 : OR2D1 port map( A1 => sec_nov_inst_m_in_l_4_port, A2 => 
                           sec_nov_inst_m_in_l_2_port, Z => 
                           sec_nov_inst_m_in_l_3_port);
   sec_nov_inst_add_239_U10 : OAI211D1 port map( A1 => 
                           sec_nov_inst_a_in_l_1_port, A2 => 
                           sec_nov_inst_a_in_r_1_port, B => 
                           sec_nov_inst_a_in_l_0_port, C => 
                           sec_nov_inst_a_in_r_0_port, Z => 
                           sec_nov_inst_add_239_n9);
   sec_nov_inst_add_239_U9 : OAI21M20D1 port map( A1 => 
                           sec_nov_inst_a_in_l_1_port, A2 => 
                           sec_nov_inst_a_in_r_1_port, B => 
                           sec_nov_inst_add_239_n9, Z => 
                           sec_nov_inst_add_239_n7);
   sec_nov_inst_add_239_U8 : OAI21D1 port map( A1 => sec_nov_inst_a_in_l_2_port
                           , A2 => sec_nov_inst_add_239_n7, B => 
                           sec_nov_inst_a_in_r_2_port, Z => 
                           sec_nov_inst_add_239_n8);
   sec_nov_inst_add_239_U7 : OAI21M20D1 port map( A1 => sec_nov_inst_add_239_n7
                           , A2 => sec_nov_inst_a_in_l_2_port, B => 
                           sec_nov_inst_add_239_n8, Z => 
                           sec_nov_inst_add_239_n5);
   sec_nov_inst_add_239_U6 : OAI21D1 port map( A1 => sec_nov_inst_a_in_l_3_port
                           , A2 => sec_nov_inst_add_239_n5, B => 
                           sec_nov_inst_a_in_r_3_port, Z => 
                           sec_nov_inst_add_239_n6);
   sec_nov_inst_add_239_U5 : OAI21M20D1 port map( A1 => sec_nov_inst_add_239_n5
                           , A2 => sec_nov_inst_a_in_l_3_port, B => 
                           sec_nov_inst_add_239_n6, Z => 
                           sec_nov_inst_add_239_n3);
   sec_nov_inst_add_239_U4 : OAI21D1 port map( A1 => sec_nov_inst_a_in_l_4_port
                           , A2 => sec_nov_inst_add_239_n3, B => 
                           sec_nov_inst_a_in_r_4_port, Z => 
                           sec_nov_inst_add_239_n4);
   sec_nov_inst_add_239_U3 : OAI21M20D1 port map( A1 => sec_nov_inst_add_239_n3
                           , A2 => sec_nov_inst_a_in_l_4_port, B => 
                           sec_nov_inst_add_239_n4, Z => 
                           sec_nov_inst_add_239_n1);
   sec_nov_inst_add_239_U2 : OAI21D1 port map( A1 => sec_nov_inst_a_in_l_5_port
                           , A2 => sec_nov_inst_add_239_n1, B => 
                           sec_nov_inst_a_in_r_5_port, Z => 
                           sec_nov_inst_add_239_n2);
   sec_nov_inst_add_239_U1 : OAI21M20D1 port map( A1 => sec_nov_inst_add_239_n1
                           , A2 => sec_nov_inst_a_in_l_5_port, B => 
                           sec_nov_inst_add_239_n2, Z => 
                           sec_nov_inst_add_239_carry_6_port);
   sec_nov_inst_add_239_U1_6 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_6_port, B => 
                           sec_nov_inst_a_in_r_6_port, CI => 
                           sec_nov_inst_add_239_carry_6_port, CO => 
                           sec_nov_inst_add_239_carry_7_port, S => 
                           sec_nov_inst_N123);
   sec_nov_inst_add_239_U1_7 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_7_port, B => 
                           sec_nov_inst_a_in_r_7_port, CI => 
                           sec_nov_inst_add_239_carry_7_port, CO => 
                           sec_nov_inst_add_239_carry_8_port, S => 
                           sec_nov_inst_N124);
   sec_nov_inst_add_239_U1_8 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_8_port, B => 
                           sec_nov_inst_a_in_r_8_port, CI => 
                           sec_nov_inst_add_239_carry_8_port, CO => 
                           sec_nov_inst_add_239_carry_9_port, S => 
                           sec_nov_inst_N125);
   sec_nov_inst_add_239_U1_9 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_9_port, B => 
                           sec_nov_inst_a_in_r_9_port, CI => 
                           sec_nov_inst_add_239_carry_9_port, CO => 
                           sec_nov_inst_add_239_carry_10_port, S => 
                           sec_nov_inst_N126);
   sec_nov_inst_add_239_U1_10 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_10_port, B => 
                           sec_nov_inst_a_in_r_10_port, CI => 
                           sec_nov_inst_add_239_carry_10_port, CO => 
                           sec_nov_inst_add_239_carry_11_port, S => 
                           sec_nov_inst_N127);
   sec_nov_inst_add_239_U1_11 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_11_port, B => 
                           sec_nov_inst_a_in_r_11_port, CI => 
                           sec_nov_inst_add_239_carry_11_port, CO => 
                           sec_nov_inst_add_239_carry_12_port, S => 
                           sec_nov_inst_N128);
   sec_nov_inst_add_239_U1_12 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_12_port, B => 
                           sec_nov_inst_a_in_r_12_port, CI => 
                           sec_nov_inst_add_239_carry_12_port, CO => 
                           sec_nov_inst_add_239_carry_13_port, S => 
                           sec_nov_inst_N129);
   sec_nov_inst_add_239_U1_13 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_13_port, B => 
                           sec_nov_inst_a_in_r_13_port, CI => 
                           sec_nov_inst_add_239_carry_13_port, CO => 
                           sec_nov_inst_add_239_carry_14_port, S => 
                           sec_nov_inst_N130);
   sec_nov_inst_add_239_U1_14 : ADFULD1 port map( A => 
                           sec_nov_inst_a_in_l_14_port, B => 
                           sec_nov_inst_a_in_r_14_port, CI => 
                           sec_nov_inst_add_239_carry_14_port, CO => 
                           sec_nov_inst_add_239_n_1009, S => sec_nov_inst_N131)
                           ;
   sec_nov_inst_mult_238_U238 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_l_6_port, A2 => 
                           sec_nov_inst_m_in_l_5_port, Z => 
                           sec_nov_inst_mult_238_n205);
   sec_nov_inst_mult_238_U237 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_7_port, A2 => 
                           sec_nov_inst_m_in_l_7_port, Z => 
                           sec_nov_inst_mult_238_n206);
   sec_nov_inst_mult_238_U236 : EXNOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_6_port, A2 => 
                           sec_nov_inst_mult_238_n201, Z => 
                           sec_nov_inst_mult_238_n241);
   sec_nov_inst_mult_238_U235 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_l_7_port, A2 => 
                           sec_nov_inst_m_in_l_6_port, Z => 
                           sec_nov_inst_mult_238_n247);
   sec_nov_inst_mult_238_U234 : NAN2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n197, A2 => 
                           sec_nov_inst_mult_238_n247, Z => 
                           sec_nov_inst_mult_238_n236);
   sec_nov_inst_mult_238_U233 : AOI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n205, A2 => 
                           sec_nov_inst_mult_238_n206, B1 => 
                           sec_nov_inst_mult_238_n241, B2 => 
                           sec_nov_inst_mult_238_n196, Z => 
                           sec_nov_inst_mult_238_n16);
   sec_nov_inst_mult_238_U232 : EXNOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_7_port, A2 => 
                           sec_nov_inst_m_in_l_5_port, Z => 
                           sec_nov_inst_mult_238_n233);
   sec_nov_inst_mult_238_U231 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_6_port, A2 => 
                           sec_nov_inst_mult_238_n195, Z => 
                           sec_nov_inst_mult_238_n232);
   sec_nov_inst_mult_238_U230 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_l_5_port, A2 => 
                           sec_nov_inst_m_in_l_4_port, Z => 
                           sec_nov_inst_mult_238_n246);
   sec_nov_inst_mult_238_U229 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n233, B1 => 
                           sec_nov_inst_mult_238_n232, B2 => 
                           sec_nov_inst_mult_238_n227, Z => 
                           sec_nov_inst_mult_238_n21);
   sec_nov_inst_mult_238_U228 : EXNOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_7_port, A2 => 
                           sec_nov_inst_m_in_l_3_port, Z => 
                           sec_nov_inst_mult_238_n223);
   sec_nov_inst_mult_238_U227 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_6_port, A2 => 
                           sec_nov_inst_mult_238_n199, Z => 
                           sec_nov_inst_mult_238_n244);
   sec_nov_inst_mult_238_U226 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_l_3_port, A2 => 
                           sec_nov_inst_m_in_l_2_port, Z => 
                           sec_nov_inst_mult_238_n245);
   sec_nov_inst_mult_238_U225 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n223, B1 => 
                           sec_nov_inst_mult_238_n244, B2 => 
                           sec_nov_inst_mult_238_n218, Z => 
                           sec_nov_inst_mult_238_n31);
   sec_nov_inst_mult_238_U224 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_2_port, A2 => 
                           sec_nov_inst_mult_238_n201, Z => 
                           sec_nov_inst_mult_238_n238);
   sec_nov_inst_mult_238_U223 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_1_port, A2 => 
                           sec_nov_inst_mult_238_n201, Z => 
                           sec_nov_inst_mult_238_n234);
   sec_nov_inst_mult_238_U222 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n197, A2 => 
                           sec_nov_inst_mult_238_n238, B1 => 
                           sec_nov_inst_mult_238_n234, B2 => 
                           sec_nov_inst_mult_238_n236, Z => 
                           sec_nov_inst_mult_238_n242);
   sec_nov_inst_mult_238_U221 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_5_port, A2 => 
                           sec_nov_inst_mult_238_n199, Z => 
                           sec_nov_inst_mult_238_n222);
   sec_nov_inst_mult_238_U220 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n244, B1 => 
                           sec_nov_inst_mult_238_n222, B2 => 
                           sec_nov_inst_mult_238_n218, Z => 
                           sec_nov_inst_mult_238_n243);
   sec_nov_inst_mult_238_U219 : OR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n242, A2 => 
                           sec_nov_inst_mult_238_n243, Z => 
                           sec_nov_inst_mult_238_n37);
   sec_nov_inst_mult_238_U218 : EXNOR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n242, A2 => 
                           sec_nov_inst_mult_238_n243, Z => 
                           sec_nov_inst_mult_238_n38);
   sec_nov_inst_mult_238_U217 : OAI32D1 port map( A1 => 
                           sec_nov_inst_mult_238_n201, A2 => 
                           sec_nov_inst_m_in_r_0_port, A3 => 
                           sec_nov_inst_mult_238_n197, B1 => 
                           sec_nov_inst_mult_238_n201, B2 => 
                           sec_nov_inst_mult_238_n236, Z => 
                           sec_nov_inst_mult_238_n57);
   sec_nov_inst_mult_238_U216 : OAI32D1 port map( A1 => 
                           sec_nov_inst_mult_238_n195, A2 => 
                           sec_nov_inst_m_in_r_0_port, A3 => 
                           sec_nov_inst_mult_238_n224, B1 => 
                           sec_nov_inst_mult_238_n195, B2 => 
                           sec_nov_inst_mult_238_n227, Z => 
                           sec_nov_inst_mult_238_n58);
   sec_nov_inst_mult_238_U215 : OAI32D1 port map( A1 => 
                           sec_nov_inst_mult_238_n199, A2 => 
                           sec_nov_inst_m_in_r_0_port, A3 => 
                           sec_nov_inst_mult_238_n215, B1 => 
                           sec_nov_inst_mult_238_n199, B2 => 
                           sec_nov_inst_mult_238_n218, Z => 
                           sec_nov_inst_mult_238_n59);
   sec_nov_inst_mult_238_U214 : OAI21D1 port map( A1 => 
                           sec_nov_inst_m_in_r_0_port, A2 => 
                           sec_nov_inst_mult_238_n202, B => 
                           sec_nov_inst_mult_238_n208, Z => 
                           sec_nov_inst_mult_238_n60);
   sec_nov_inst_mult_238_U213 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_5_port, A2 => 
                           sec_nov_inst_mult_238_n201, Z => 
                           sec_nov_inst_mult_238_n240);
   sec_nov_inst_mult_238_U212 : OAI22M10D1 port map( A1 => 
                           sec_nov_inst_mult_238_n241, A2 => 
                           sec_nov_inst_mult_238_n197, B1 => 
                           sec_nov_inst_mult_238_n240, B2 => 
                           sec_nov_inst_mult_238_n236, Z => 
                           sec_nov_inst_mult_238_n62);
   sec_nov_inst_mult_238_U211 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_4_port, A2 => 
                           sec_nov_inst_mult_238_n201, Z => 
                           sec_nov_inst_mult_238_n239);
   sec_nov_inst_mult_238_U210 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n197, A2 => 
                           sec_nov_inst_mult_238_n240, B1 => 
                           sec_nov_inst_mult_238_n239, B2 => 
                           sec_nov_inst_mult_238_n236, Z => 
                           sec_nov_inst_mult_238_n63);
   sec_nov_inst_mult_238_U209 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_3_port, A2 => 
                           sec_nov_inst_mult_238_n201, Z => 
                           sec_nov_inst_mult_238_n237);
   sec_nov_inst_mult_238_U208 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n197, A2 => 
                           sec_nov_inst_mult_238_n239, B1 => 
                           sec_nov_inst_mult_238_n237, B2 => 
                           sec_nov_inst_mult_238_n236, Z => 
                           sec_nov_inst_mult_238_n64);
   sec_nov_inst_mult_238_U207 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n197, A2 => 
                           sec_nov_inst_mult_238_n237, B1 => 
                           sec_nov_inst_mult_238_n238, B2 => 
                           sec_nov_inst_mult_238_n236, Z => 
                           sec_nov_inst_mult_238_n65);
   sec_nov_inst_mult_238_U206 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n201, A2 => 
                           sec_nov_inst_m_in_r_0_port, Z => 
                           sec_nov_inst_mult_238_n235);
   sec_nov_inst_mult_238_U205 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n197, A2 => 
                           sec_nov_inst_mult_238_n234, B1 => 
                           sec_nov_inst_mult_238_n235, B2 => 
                           sec_nov_inst_mult_238_n236, Z => 
                           sec_nov_inst_mult_238_n67);
   sec_nov_inst_mult_238_U204 : NOR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n197, A2 => 
                           sec_nov_inst_mult_238_n203, Z => 
                           sec_nov_inst_mult_238_n68);
   sec_nov_inst_mult_238_U203 : AO21D1 port map( A1 => 
                           sec_nov_inst_mult_238_n227, A2 => 
                           sec_nov_inst_mult_238_n224, B => 
                           sec_nov_inst_mult_238_n233, Z => 
                           sec_nov_inst_mult_238_n69);
   sec_nov_inst_mult_238_U202 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_5_port, A2 => 
                           sec_nov_inst_mult_238_n195, Z => 
                           sec_nov_inst_mult_238_n231);
   sec_nov_inst_mult_238_U201 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n232, B1 => 
                           sec_nov_inst_mult_238_n231, B2 => 
                           sec_nov_inst_mult_238_n227, Z => 
                           sec_nov_inst_mult_238_n70);
   sec_nov_inst_mult_238_U200 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_4_port, A2 => 
                           sec_nov_inst_mult_238_n195, Z => 
                           sec_nov_inst_mult_238_n230);
   sec_nov_inst_mult_238_U199 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n231, B1 => 
                           sec_nov_inst_mult_238_n230, B2 => 
                           sec_nov_inst_mult_238_n227, Z => 
                           sec_nov_inst_mult_238_n71);
   sec_nov_inst_mult_238_U198 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_3_port, A2 => 
                           sec_nov_inst_mult_238_n195, Z => 
                           sec_nov_inst_mult_238_n229);
   sec_nov_inst_mult_238_U197 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n230, B1 => 
                           sec_nov_inst_mult_238_n229, B2 => 
                           sec_nov_inst_mult_238_n227, Z => 
                           sec_nov_inst_mult_238_n72);
   sec_nov_inst_mult_238_U196 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_2_port, A2 => 
                           sec_nov_inst_mult_238_n195, Z => 
                           sec_nov_inst_mult_238_n228);
   sec_nov_inst_mult_238_U195 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n229, B1 => 
                           sec_nov_inst_mult_238_n228, B2 => 
                           sec_nov_inst_mult_238_n227, Z => 
                           sec_nov_inst_mult_238_n73);
   sec_nov_inst_mult_238_U194 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_1_port, A2 => 
                           sec_nov_inst_mult_238_n195, Z => 
                           sec_nov_inst_mult_238_n225);
   sec_nov_inst_mult_238_U193 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n228, B1 => 
                           sec_nov_inst_mult_238_n225, B2 => 
                           sec_nov_inst_mult_238_n227, Z => 
                           sec_nov_inst_mult_238_n74);
   sec_nov_inst_mult_238_U192 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n195, A2 => 
                           sec_nov_inst_m_in_r_0_port, Z => 
                           sec_nov_inst_mult_238_n226);
   sec_nov_inst_mult_238_U191 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n225, B1 => 
                           sec_nov_inst_mult_238_n226, B2 => 
                           sec_nov_inst_mult_238_n227, Z => 
                           sec_nov_inst_mult_238_n75);
   sec_nov_inst_mult_238_U190 : NOR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n203, Z => 
                           sec_nov_inst_mult_238_n76);
   sec_nov_inst_mult_238_U189 : AO21D1 port map( A1 => 
                           sec_nov_inst_mult_238_n218, A2 => 
                           sec_nov_inst_mult_238_n215, B => 
                           sec_nov_inst_mult_238_n223, Z => 
                           sec_nov_inst_mult_238_n77);
   sec_nov_inst_mult_238_U188 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_4_port, A2 => 
                           sec_nov_inst_mult_238_n199, Z => 
                           sec_nov_inst_mult_238_n221);
   sec_nov_inst_mult_238_U187 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n222, B1 => 
                           sec_nov_inst_mult_238_n221, B2 => 
                           sec_nov_inst_mult_238_n218, Z => 
                           sec_nov_inst_mult_238_n79);
   sec_nov_inst_mult_238_U186 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_3_port, A2 => 
                           sec_nov_inst_mult_238_n199, Z => 
                           sec_nov_inst_mult_238_n220);
   sec_nov_inst_mult_238_U185 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n221, B1 => 
                           sec_nov_inst_mult_238_n220, B2 => 
                           sec_nov_inst_mult_238_n218, Z => 
                           sec_nov_inst_mult_238_n80);
   sec_nov_inst_mult_238_U184 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_2_port, A2 => 
                           sec_nov_inst_mult_238_n199, Z => 
                           sec_nov_inst_mult_238_n219);
   sec_nov_inst_mult_238_U183 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n220, B1 => 
                           sec_nov_inst_mult_238_n219, B2 => 
                           sec_nov_inst_mult_238_n218, Z => 
                           sec_nov_inst_mult_238_n81);
   sec_nov_inst_mult_238_U182 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_1_port, A2 => 
                           sec_nov_inst_mult_238_n199, Z => 
                           sec_nov_inst_mult_238_n216);
   sec_nov_inst_mult_238_U181 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n219, B1 => 
                           sec_nov_inst_mult_238_n216, B2 => 
                           sec_nov_inst_mult_238_n218, Z => 
                           sec_nov_inst_mult_238_n82);
   sec_nov_inst_mult_238_U180 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n199, A2 => 
                           sec_nov_inst_m_in_r_0_port, Z => 
                           sec_nov_inst_mult_238_n217);
   sec_nov_inst_mult_238_U179 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n216, B1 => 
                           sec_nov_inst_mult_238_n217, B2 => 
                           sec_nov_inst_mult_238_n218, Z => 
                           sec_nov_inst_mult_238_n83);
   sec_nov_inst_mult_238_U178 : NOR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n203, Z => 
                           sec_nov_inst_mult_238_n84);
   sec_nov_inst_mult_238_U177 : EXNOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_7_port, A2 => 
                           sec_nov_inst_m_in_l_1_port, Z => 
                           sec_nov_inst_mult_238_n214);
   sec_nov_inst_mult_238_U176 : AO21D1 port map( A1 => 
                           sec_nov_inst_mult_238_n200, A2 => 
                           sec_nov_inst_mult_238_n208, B => 
                           sec_nov_inst_mult_238_n214, Z => 
                           sec_nov_inst_mult_238_n85);
   sec_nov_inst_mult_238_U175 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_6_port, A2 => 
                           sec_nov_inst_mult_238_n202, Z => 
                           sec_nov_inst_mult_238_n213);
   sec_nov_inst_mult_238_U174 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n214, A2 => 
                           sec_nov_inst_mult_238_n200, B1 => 
                           sec_nov_inst_mult_238_n213, B2 => 
                           sec_nov_inst_mult_238_n208, Z => 
                           sec_nov_inst_mult_238_n86);
   sec_nov_inst_mult_238_U173 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_5_port, A2 => 
                           sec_nov_inst_mult_238_n202, Z => 
                           sec_nov_inst_mult_238_n212);
   sec_nov_inst_mult_238_U172 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n213, A2 => 
                           sec_nov_inst_mult_238_n200, B1 => 
                           sec_nov_inst_mult_238_n212, B2 => 
                           sec_nov_inst_mult_238_n208, Z => 
                           sec_nov_inst_mult_238_n87);
   sec_nov_inst_mult_238_U171 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_4_port, A2 => 
                           sec_nov_inst_mult_238_n202, Z => 
                           sec_nov_inst_mult_238_n211);
   sec_nov_inst_mult_238_U170 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n212, A2 => 
                           sec_nov_inst_mult_238_n200, B1 => 
                           sec_nov_inst_mult_238_n211, B2 => 
                           sec_nov_inst_mult_238_n208, Z => 
                           sec_nov_inst_mult_238_n88);
   sec_nov_inst_mult_238_U169 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_3_port, A2 => 
                           sec_nov_inst_mult_238_n202, Z => 
                           sec_nov_inst_mult_238_n210);
   sec_nov_inst_mult_238_U168 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n211, A2 => 
                           sec_nov_inst_mult_238_n200, B1 => 
                           sec_nov_inst_mult_238_n210, B2 => 
                           sec_nov_inst_mult_238_n208, Z => 
                           sec_nov_inst_mult_238_n89);
   sec_nov_inst_mult_238_U167 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_2_port, A2 => 
                           sec_nov_inst_mult_238_n202, Z => 
                           sec_nov_inst_mult_238_n209);
   sec_nov_inst_mult_238_U166 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n210, A2 => 
                           sec_nov_inst_mult_238_n200, B1 => 
                           sec_nov_inst_mult_238_n209, B2 => 
                           sec_nov_inst_mult_238_n208, Z => 
                           sec_nov_inst_mult_238_n90);
   sec_nov_inst_mult_238_U165 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_r_1_port, A2 => 
                           sec_nov_inst_mult_238_n202, Z => 
                           sec_nov_inst_mult_238_n207);
   sec_nov_inst_mult_238_U164 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n209, A2 => 
                           sec_nov_inst_mult_238_n200, B1 => 
                           sec_nov_inst_mult_238_n207, B2 => 
                           sec_nov_inst_mult_238_n208, Z => 
                           sec_nov_inst_mult_238_n91);
   sec_nov_inst_mult_238_U163 : OAI22D1 port map( A1 => 
                           sec_nov_inst_mult_238_n207, A2 => 
                           sec_nov_inst_mult_238_n200, B1 => 
                           sec_nov_inst_m_in_r_0_port, B2 => 
                           sec_nov_inst_mult_238_n208, Z => 
                           sec_nov_inst_mult_238_n92);
   sec_nov_inst_mult_238_U162 : NOR2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n200, A2 => 
                           sec_nov_inst_mult_238_n203, Z => 
                           sec_nov_inst_m_out_0_port);
   sec_nov_inst_mult_238_U161 : OAI21D1 port map( A1 => 
                           sec_nov_inst_mult_238_n196, A2 => 
                           sec_nov_inst_mult_238_n205, B => 
                           sec_nov_inst_mult_238_n206, Z => 
                           sec_nov_inst_mult_238_n204);
   sec_nov_inst_mult_238_U160 : EXNOR3D1 port map( A1 => 
                           sec_nov_inst_mult_238_n2, A2 => 
                           sec_nov_inst_mult_238_n16, A3 => 
                           sec_nov_inst_mult_238_n204, Z => 
                           sec_nov_inst_m_out_14_port);
   sec_nov_inst_mult_238_U159 : INVD1 port map( A => sec_nov_inst_m_in_r_0_port
                           , Z => sec_nov_inst_mult_238_n203);
   sec_nov_inst_mult_238_U158 : INVD1 port map( A => sec_nov_inst_mult_238_n21,
                           Z => sec_nov_inst_mult_238_n194);
   sec_nov_inst_mult_238_U157 : INVD1 port map( A => sec_nov_inst_mult_238_n31,
                           Z => sec_nov_inst_mult_238_n198);
   sec_nov_inst_mult_238_U156 : NAN2D1 port map( A1 => 
                           sec_nov_inst_m_in_l_1_port, A2 => 
                           sec_nov_inst_mult_238_n200, Z => 
                           sec_nov_inst_mult_238_n208);
   sec_nov_inst_mult_238_U155 : INVD1 port map( A => sec_nov_inst_m_in_l_1_port
                           , Z => sec_nov_inst_mult_238_n202);
   sec_nov_inst_mult_238_U154 : INVD1 port map( A => sec_nov_inst_mult_238_n236
                           , Z => sec_nov_inst_mult_238_n196);
   sec_nov_inst_mult_238_U153 : INVD1 port map( A => sec_nov_inst_m_in_l_7_port
                           , Z => sec_nov_inst_mult_238_n201);
   sec_nov_inst_mult_238_U152 : INVD1 port map( A => sec_nov_inst_m_in_l_5_port
                           , Z => sec_nov_inst_mult_238_n195);
   sec_nov_inst_mult_238_U151 : INVD1 port map( A => sec_nov_inst_mult_238_n205
                           , Z => sec_nov_inst_mult_238_n197);
   sec_nov_inst_mult_238_U150 : INVD1 port map( A => sec_nov_inst_m_in_l_0_port
                           , Z => sec_nov_inst_mult_238_n200);
   sec_nov_inst_mult_238_U149 : NAN2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n215, A2 => 
                           sec_nov_inst_mult_238_n245, Z => 
                           sec_nov_inst_mult_238_n218);
   sec_nov_inst_mult_238_U148 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_l_2_port, A2 => 
                           sec_nov_inst_mult_238_n202, Z => 
                           sec_nov_inst_mult_238_n215);
   sec_nov_inst_mult_238_U147 : NAN2D1 port map( A1 => 
                           sec_nov_inst_mult_238_n224, A2 => 
                           sec_nov_inst_mult_238_n246, Z => 
                           sec_nov_inst_mult_238_n227);
   sec_nov_inst_mult_238_U146 : EXOR2D1 port map( A1 => 
                           sec_nov_inst_m_in_l_4_port, A2 => 
                           sec_nov_inst_mult_238_n199, Z => 
                           sec_nov_inst_mult_238_n224);
   sec_nov_inst_mult_238_U145 : INVD1 port map( A => sec_nov_inst_m_in_l_3_port
                           , Z => sec_nov_inst_mult_238_n199);
   sec_nov_inst_mult_238_U37 : ADHALFDL port map( A => 
                           sec_nov_inst_mult_238_n83, B => 
                           sec_nov_inst_mult_238_n90, CO => 
                           sec_nov_inst_mult_238_n55, S => 
                           sec_nov_inst_mult_238_n56);
   sec_nov_inst_mult_238_U36 : ADFULD1 port map( A => sec_nov_inst_mult_238_n89
                           , B => sec_nov_inst_mult_238_n76, CI => 
                           sec_nov_inst_mult_238_n82, CO => 
                           sec_nov_inst_mult_238_n53, S => 
                           sec_nov_inst_mult_238_n54);
   sec_nov_inst_mult_238_U35 : ADHALFDL port map( A => 
                           sec_nov_inst_mult_238_n58, B => 
                           sec_nov_inst_mult_238_n88, CO => 
                           sec_nov_inst_mult_238_n51, S => 
                           sec_nov_inst_mult_238_n52);
   sec_nov_inst_mult_238_U34 : ADFULD1 port map( A => sec_nov_inst_mult_238_n75
                           , B => sec_nov_inst_mult_238_n81, CI => 
                           sec_nov_inst_mult_238_n52, CO => 
                           sec_nov_inst_mult_238_n49, S => 
                           sec_nov_inst_mult_238_n50);
   sec_nov_inst_mult_238_U33 : ADFULD1 port map( A => sec_nov_inst_mult_238_n87
                           , B => sec_nov_inst_mult_238_n68, CI => 
                           sec_nov_inst_mult_238_n80, CO => 
                           sec_nov_inst_mult_238_n47, S => 
                           sec_nov_inst_mult_238_n48);
   sec_nov_inst_mult_238_U32 : ADFULD1 port map( A => sec_nov_inst_mult_238_n51
                           , B => sec_nov_inst_mult_238_n74, CI => 
                           sec_nov_inst_mult_238_n48, CO => 
                           sec_nov_inst_mult_238_n45, S => 
                           sec_nov_inst_mult_238_n46);
   sec_nov_inst_mult_238_U31 : ADHALFDL port map( A => 
                           sec_nov_inst_mult_238_n57, B => 
                           sec_nov_inst_mult_238_n86, CO => 
                           sec_nov_inst_mult_238_n43, S => 
                           sec_nov_inst_mult_238_n44);
   sec_nov_inst_mult_238_U30 : ADFULD1 port map( A => sec_nov_inst_mult_238_n67
                           , B => sec_nov_inst_mult_238_n79, CI => 
                           sec_nov_inst_mult_238_n73, CO => 
                           sec_nov_inst_mult_238_n41, S => 
                           sec_nov_inst_mult_238_n42);
   sec_nov_inst_mult_238_U29 : ADFULD1 port map( A => sec_nov_inst_mult_238_n47
                           , B => sec_nov_inst_mult_238_n44, CI => 
                           sec_nov_inst_mult_238_n42, CO => 
                           sec_nov_inst_mult_238_n39, S => 
                           sec_nov_inst_mult_238_n40);
   sec_nov_inst_mult_238_U26 : ADFULD1 port map( A => sec_nov_inst_mult_238_n85
                           , B => sec_nov_inst_mult_238_n72, CI => 
                           sec_nov_inst_mult_238_n43, CO => 
                           sec_nov_inst_mult_238_n35, S => 
                           sec_nov_inst_mult_238_n36);
   sec_nov_inst_mult_238_U25 : ADFULD1 port map( A => sec_nov_inst_mult_238_n41
                           , B => sec_nov_inst_mult_238_n38, CI => 
                           sec_nov_inst_mult_238_n36, CO => 
                           sec_nov_inst_mult_238_n33, S => 
                           sec_nov_inst_mult_238_n34);
   sec_nov_inst_mult_238_U23 : ADFULD1 port map( A => sec_nov_inst_mult_238_n65
                           , B => sec_nov_inst_mult_238_n71, CI => 
                           sec_nov_inst_mult_238_n198, CO => 
                           sec_nov_inst_mult_238_n29, S => 
                           sec_nov_inst_mult_238_n30);
   sec_nov_inst_mult_238_U22 : ADFULD1 port map( A => sec_nov_inst_mult_238_n35
                           , B => sec_nov_inst_mult_238_n37, CI => 
                           sec_nov_inst_mult_238_n30, CO => 
                           sec_nov_inst_mult_238_n27, S => 
                           sec_nov_inst_mult_238_n28);
   sec_nov_inst_mult_238_U21 : ADFULD1 port map( A => sec_nov_inst_mult_238_n70
                           , B => sec_nov_inst_mult_238_n31, CI => 
                           sec_nov_inst_mult_238_n64, CO => 
                           sec_nov_inst_mult_238_n25, S => 
                           sec_nov_inst_mult_238_n26);
   sec_nov_inst_mult_238_U20 : ADFULD1 port map( A => sec_nov_inst_mult_238_n29
                           , B => sec_nov_inst_mult_238_n77, CI => 
                           sec_nov_inst_mult_238_n26, CO => 
                           sec_nov_inst_mult_238_n23, S => 
                           sec_nov_inst_mult_238_n24);
   sec_nov_inst_mult_238_U18 : ADFULD1 port map( A => 
                           sec_nov_inst_mult_238_n194, B => 
                           sec_nov_inst_mult_238_n63, CI => 
                           sec_nov_inst_mult_238_n25, CO => 
                           sec_nov_inst_mult_238_n19, S => 
                           sec_nov_inst_mult_238_n20);
   sec_nov_inst_mult_238_U17 : ADFULD1 port map( A => sec_nov_inst_mult_238_n62
                           , B => sec_nov_inst_mult_238_n21, CI => 
                           sec_nov_inst_mult_238_n69, CO => 
                           sec_nov_inst_mult_238_n17, S => 
                           sec_nov_inst_mult_238_n18);
   sec_nov_inst_mult_238_U15 : ADHALFDL port map( A => 
                           sec_nov_inst_mult_238_n92, B => 
                           sec_nov_inst_mult_238_n60, CO => 
                           sec_nov_inst_mult_238_n14, S => 
                           sec_nov_inst_m_out_1_port);
   sec_nov_inst_mult_238_U14 : ADFULD1 port map( A => sec_nov_inst_mult_238_n91
                           , B => sec_nov_inst_mult_238_n84, CI => 
                           sec_nov_inst_mult_238_n14, CO => 
                           sec_nov_inst_mult_238_n13, S => 
                           sec_nov_inst_m_out_2_port);
   sec_nov_inst_mult_238_U13 : ADFULD1 port map( A => sec_nov_inst_mult_238_n56
                           , B => sec_nov_inst_mult_238_n59, CI => 
                           sec_nov_inst_mult_238_n13, CO => 
                           sec_nov_inst_mult_238_n12, S => 
                           sec_nov_inst_m_out_3_port);
   sec_nov_inst_mult_238_U12 : ADFULD1 port map( A => sec_nov_inst_mult_238_n54
                           , B => sec_nov_inst_mult_238_n55, CI => 
                           sec_nov_inst_mult_238_n12, CO => 
                           sec_nov_inst_mult_238_n11, S => 
                           sec_nov_inst_m_out_4_port);
   sec_nov_inst_mult_238_U11 : ADFULD1 port map( A => sec_nov_inst_mult_238_n50
                           , B => sec_nov_inst_mult_238_n53, CI => 
                           sec_nov_inst_mult_238_n11, CO => 
                           sec_nov_inst_mult_238_n10, S => 
                           sec_nov_inst_m_out_5_port);
   sec_nov_inst_mult_238_U10 : ADFULD1 port map( A => sec_nov_inst_mult_238_n46
                           , B => sec_nov_inst_mult_238_n49, CI => 
                           sec_nov_inst_mult_238_n10, CO => 
                           sec_nov_inst_mult_238_n9, S => 
                           sec_nov_inst_m_out_6_port);
   sec_nov_inst_mult_238_U9 : ADFULD1 port map( A => sec_nov_inst_mult_238_n40,
                           B => sec_nov_inst_mult_238_n45, CI => 
                           sec_nov_inst_mult_238_n9, CO => 
                           sec_nov_inst_mult_238_n8, S => 
                           sec_nov_inst_m_out_7_port);
   sec_nov_inst_mult_238_U8 : ADFULD1 port map( A => sec_nov_inst_mult_238_n34,
                           B => sec_nov_inst_mult_238_n39, CI => 
                           sec_nov_inst_mult_238_n8, CO => 
                           sec_nov_inst_mult_238_n7, S => 
                           sec_nov_inst_m_out_8_port);
   sec_nov_inst_mult_238_U7 : ADFULD1 port map( A => sec_nov_inst_mult_238_n28,
                           B => sec_nov_inst_mult_238_n33, CI => 
                           sec_nov_inst_mult_238_n7, CO => 
                           sec_nov_inst_mult_238_n6, S => 
                           sec_nov_inst_m_out_9_port);
   sec_nov_inst_mult_238_U6 : ADFULD1 port map( A => sec_nov_inst_mult_238_n24,
                           B => sec_nov_inst_mult_238_n27, CI => 
                           sec_nov_inst_mult_238_n6, CO => 
                           sec_nov_inst_mult_238_n5, S => 
                           sec_nov_inst_m_out_10_port);
   sec_nov_inst_mult_238_U5 : ADFULD1 port map( A => sec_nov_inst_mult_238_n20,
                           B => sec_nov_inst_mult_238_n23, CI => 
                           sec_nov_inst_mult_238_n5, CO => 
                           sec_nov_inst_mult_238_n4, S => 
                           sec_nov_inst_m_out_11_port);
   sec_nov_inst_mult_238_U4 : ADFULD1 port map( A => sec_nov_inst_mult_238_n19,
                           B => sec_nov_inst_mult_238_n18, CI => 
                           sec_nov_inst_mult_238_n4, CO => 
                           sec_nov_inst_mult_238_n3, S => 
                           sec_nov_inst_m_out_12_port);
   sec_nov_inst_mult_238_U3 : ADFULD1 port map( A => sec_nov_inst_mult_238_n17,
                           B => sec_nov_inst_mult_238_n16, CI => 
                           sec_nov_inst_mult_238_n3, CO => 
                           sec_nov_inst_mult_238_n2, S => 
                           sec_nov_inst_m_out_13_port);

end flat_rtl_none_10;
