
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_TRA3 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type SIGNED is array (INTEGER range <>) of std_logic;

end CONV_PACK_TRA3;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture flat_rtl_none_10 of TRA3 is

   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVBD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal arx_i1_reg_7_port, arx_i1_reg_6_port, arx_i1_reg_5_port, 
      arx_i1_reg_4_port, arx_i1_reg_3_port, arx_i1_reg_2_port, 
      arx_i1_reg_1_port, arx_i1_reg_0_port, arx_r1_reg_14_port, 
      arx_r1_reg_13_port, arx_r1_reg_12_port, arx_r1_reg_11_port, 
      arx_r1_reg_10_port, arx_r1_reg_9_port, arx_r1_reg_8_port, 
      arx_r1_reg_7_port, arx_r1_reg_6_port, arx_r1_reg_5_port, 
      arx_r1_reg_4_port, arx_r1_reg_3_port, arx_r1_reg_2_port, 
      arx_r1_reg_1_port, arx_r1_reg_0_port, arx_r2_reg_14_port, 
      arx_r2_reg_13_port, arx_r2_reg_12_port, arx_r2_reg_11_port, 
      arx_r2_reg_10_port, arx_r2_reg_9_port, arx_r2_reg_8_port, 
      arx_r2_reg_7_port, arx_r2_reg_6_port, arx_r2_reg_5_port, 
      arx_r2_reg_4_port, arx_r2_reg_3_port, arx_r2_reg_2_port, 
      arx_r2_reg_1_port, arx_r2_reg_0_port, arx_r3_reg_14_port, 
      arx_r3_reg_13_port, arx_r3_reg_12_port, arx_r3_reg_11_port, 
      arx_r3_reg_10_port, arx_r3_reg_9_port, arx_r3_reg_8_port, 
      arx_r3_reg_7_port, arx_r3_reg_6_port, arx_r3_reg_5_port, 
      arx_r3_reg_4_port, arx_r3_reg_3_port, arx_r3_reg_2_port, 
      arx_r3_reg_1_port, arx_r3_reg_0_port, arx_r4_reg_14_port, 
      arx_r4_reg_13_port, arx_r4_reg_12_port, arx_r4_reg_11_port, 
      arx_r4_reg_10_port, arx_r4_reg_9_port, arx_r4_reg_8_port, 
      arx_r4_reg_7_port, arx_r4_reg_6_port, arx_r4_reg_5_port, 
      arx_r4_reg_4_port, arx_r4_reg_3_port, arx_r4_reg_2_port, 
      arx_r4_reg_1_port, arx_d1_reg_14_port, arx_d1_reg_13_port, 
      arx_d1_reg_12_port, arx_d1_reg_11_port, arx_d1_reg_10_port, 
      arx_d1_reg_9_port, arx_d1_reg_8_port, arx_d1_reg_7_port, 
      arx_d2_reg_14_port, arx_d2_reg_13_port, arx_d2_reg_12_port, 
      arx_d2_reg_11_port, arx_d2_reg_10_port, arx_d2_reg_9_port, 
      arx_d2_reg_8_port, arx_d2_reg_7_port, arx_state_reg_1_port, 
      arx_state_reg_0_port, m1_in_r_7_port, m1_in_r_6_port, m1_in_r_5_port, 
      m1_in_r_4_port, m1_in_r_3_port, m1_in_r_2_port, m1_in_r_1_port, 
      m1_in_r_0_port, m1_out_15, m1_out_12_port, m1_out_11_port, m1_out_10_port
      , m1_out_9_port, m1_out_8_port, m1_out_7_port, m1_out_6_port, 
      m1_out_5_port, m1_out_4_port, m1_out_3_port, m1_out_2_port, m1_out_1_port
      , m1_out_0_port, m2_in_r_7_port, m2_in_r_6_port, m2_in_r_5_port, 
      m2_in_r_4_port, m2_in_r_3_port, m2_in_r_2_port, m2_in_r_1_port, 
      m2_in_r_0_port, m2_out_14_port, m2_out_13_port, m2_out_12_port, 
      m2_out_11_port, m2_out_10_port, m2_out_9_port, m2_out_8_port, 
      m2_out_7_port, m2_out_6_port, m2_out_5_port, m2_out_4_port, m2_out_3_port
      , m2_out_2_port, m2_out_1_port, m2_out_0_port, m3_out_14_port, 
      m3_out_13_port, m3_out_12_port, m3_out_11_port, m3_out_10_port, 
      m3_out_9_port, m3_out_8_port, m3_out_7_port, m3_out_6_port, m3_out_5_port
      , m3_out_4_port, m3_out_3_port, m3_out_2_port, m3_out_1_port, 
      m4_in_r_7_port, m4_in_r_6_port, m4_in_r_5_port, m4_in_r_4_port, 
      m4_in_r_3_port, m4_in_r_2_port, m4_in_r_1_port, m4_in_r_0_port, 
      m4_out_14_port, m4_out_13_port, m4_out_12_port, m4_out_11_port, 
      m4_out_10_port, m4_out_9_port, m4_out_8_port, m4_out_7_port, 
      m4_out_6_port, m4_out_5_port, m4_out_4_port, m4_out_3_port, m4_out_2_port
      , m4_out_1_port, m4_out_0_port, m5_in_l_0, m5_in_r_7_port, m5_in_r_6_port
      , m5_in_r_5_port, m5_in_r_4_port, m5_in_r_3_port, m5_in_r_2_port, 
      m5_in_r_1_port, m5_in_r_0_port, m5_out_15, m5_out_12_port, m5_out_11_port
      , m5_out_10_port, m5_out_9_port, m5_out_8_port, m5_out_7_port, 
      m5_out_6_port, m5_out_5_port, m5_out_4_port, m5_out_3_port, m5_out_2_port
      , m5_out_1_port, m5_out_0_port, a1_in_l_14_port, a1_in_l_13_port, 
      a1_in_l_12_port, a1_in_l_11_port, a1_in_l_10_port, a1_in_l_9_port, 
      a1_in_l_8_port, a1_in_l_7_port, a1_in_l_6_port, a1_in_l_5_port, 
      a1_in_l_4_port, a1_in_l_3_port, a1_in_l_2_port, a1_in_l_1_port, 
      a1_in_l_0_port, a1_in_r_14_port, a1_in_r_13_port, a1_in_r_12_port, 
      a1_in_r_11_port, a1_in_r_10_port, a1_in_r_9_port, a1_in_r_8_port, 
      a1_in_r_7_port, a1_in_r_6_port, a1_in_r_5_port, a1_in_r_4_port, 
      a1_in_r_3_port, a1_in_r_2_port, a1_in_r_1_port, a1_in_r_0_port, 
      a1_out_7_port, a1_out_6_port, a1_out_5_port, a1_out_4_port, a1_out_3_port
      , a1_out_2_port, a1_out_1_port, a1_out_0_port, a2_in_l_14_port, 
      a2_in_l_13_port, a2_in_l_12_port, a2_in_l_11_port, a2_in_l_10_port, 
      a2_in_l_9_port, a2_in_l_8_port, a2_in_l_7_port, a2_in_l_6_port, 
      a2_in_l_5_port, a2_in_l_4_port, a2_in_l_3_port, a2_in_l_2_port, 
      a2_in_l_1_port, a2_in_l_0_port, a2_in_r_14_port, a2_in_r_13_port, 
      a2_in_r_12_port, a2_in_r_11_port, a2_in_r_10_port, a2_in_r_9_port, 
      a2_in_r_8_port, a2_in_r_7_port, a2_in_r_6_port, a2_in_r_5_port, 
      a2_in_r_4_port, a2_in_r_3_port, a2_in_r_2_port, a2_in_r_1_port, 
      a2_in_r_0_port, a2_out_7_port, a2_out_6_port, a2_out_5_port, 
      a2_out_4_port, a2_out_3_port, a2_out_2_port, a2_out_1_port, a2_out_0_port
      , state_0, N44, N45, N46, N47, N48, N49, N50, N51, N106, N107, N108, N109
      , N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
      N122, N123, net1801, n92, n94, n95, n96, n97, n98, n99, n100, n101, n102,
      n103, n104, n105, n1060, n1070, n1080, n1090, n1100, n1110, n1120, n1130,
      n1140, n1150, n1160, n1170, n1180, n1190, n1200, n1210, n1220, n1230, 
      n124, n125, n126, n127, n129, n130, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, add_416_C244_rn_carry_1_port, 
      add_416_C244_rn_carry_2_port, add_416_C244_rn_carry_3_port, 
      add_416_C244_rn_carry_4_port, add_416_C244_rn_carry_5_port, 
      add_416_C244_rn_carry_6_port, add_416_C244_rn_carry_7_port, 
      add_416_C243_rn_carry_1_port, add_416_C243_rn_carry_2_port, 
      add_416_C243_rn_carry_3_port, add_416_C243_rn_carry_4_port, 
      add_416_C243_rn_carry_5_port, add_416_C243_rn_carry_6_port, 
      add_416_C243_rn_carry_7_port, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n_1037, n_1038, n_1039, n_1040, n_1041, 
      n_1042, n_1043, n_1044, n_1045, n_1046, n_1047, n_1048, n_1049, n_1050, 
      n_1051, n_1052, n_1053, n_1054, add_244_n9, add_244_n8, add_244_n7, 
      add_244_n6, add_244_n5, add_244_n4, add_244_n3, add_244_n2, add_244_n1, 
      add_244_carry_6_port, add_244_carry_7_port, add_244_carry_8_port, 
      add_244_carry_9_port, add_244_carry_10_port, add_244_carry_11_port, 
      add_244_carry_12_port, add_244_carry_13_port, add_244_carry_14_port, 
      add_243_n9, add_243_n8, add_243_n7, add_243_n6, add_243_n5, add_243_n4, 
      add_243_n3, add_243_n2, add_243_n1, add_243_carry_6_port, 
      add_243_carry_7_port, add_243_carry_8_port, add_243_carry_9_port, 
      add_243_carry_10_port, add_243_carry_11_port, add_243_carry_12_port, 
      add_243_carry_13_port, add_243_carry_14_port, mult_238_n130, 
      mult_238_n129, mult_238_n128, mult_238_n127, mult_238_n126, mult_238_n125
      , mult_238_n124, mult_238_n123, mult_238_n122, mult_238_n121, 
      mult_238_n119, mult_238_n71, mult_238_n70, mult_238_n69, mult_238_n68, 
      mult_238_n67, mult_238_n66, mult_238_n65, mult_238_n64, mult_238_n63, 
      mult_238_n62, mult_238_n61, mult_238_n60, mult_238_n59, mult_238_n58, 
      mult_238_n57, mult_238_n56, mult_238_n55, mult_238_n54, mult_238_n53, 
      mult_238_n52, mult_238_n51, mult_238_n50, mult_238_n49, mult_238_n48, 
      mult_238_n47, mult_238_n46, mult_238_n45, mult_238_n44, mult_238_n43, 
      mult_238_n42, mult_238_n41, mult_238_n40, mult_238_n39, mult_238_n38, 
      mult_238_n37, mult_238_n36, mult_238_n35, mult_238_n33, mult_238_n32, 
      mult_238_n31, mult_238_n30, mult_238_n29, mult_238_n27, mult_238_n26, 
      mult_238_n25, mult_238_n24, mult_238_n23, mult_238_n21, mult_238_n20, 
      mult_238_n19, mult_238_n18, mult_238_n17, mult_238_n16, mult_238_n15, 
      mult_238_n14, mult_238_n13, mult_238_n12, mult_238_n11, mult_238_n10, 
      mult_238_n9, mult_238_n8, mult_238_n7, mult_238_n6, mult_238_n5, 
      mult_238_n4, mult_238_n3, mult_238_n2, mult_242_n130, mult_242_n129, 
      mult_242_n128, mult_242_n127, mult_242_n126, mult_242_n125, mult_242_n124
      , mult_242_n123, mult_242_n122, mult_242_n121, mult_242_n119, 
      mult_242_n71, mult_242_n70, mult_242_n69, mult_242_n68, mult_242_n67, 
      mult_242_n66, mult_242_n65, mult_242_n64, mult_242_n63, mult_242_n62, 
      mult_242_n61, mult_242_n60, mult_242_n59, mult_242_n58, mult_242_n57, 
      mult_242_n56, mult_242_n55, mult_242_n54, mult_242_n53, mult_242_n52, 
      mult_242_n51, mult_242_n50, mult_242_n49, mult_242_n48, mult_242_n47, 
      mult_242_n46, mult_242_n45, mult_242_n44, mult_242_n43, mult_242_n42, 
      mult_242_n41, mult_242_n40, mult_242_n39, mult_242_n38, mult_242_n37, 
      mult_242_n36, mult_242_n35, mult_242_n33, mult_242_n32, mult_242_n31, 
      mult_242_n30, mult_242_n29, mult_242_n27, mult_242_n26, mult_242_n25, 
      mult_242_n24, mult_242_n23, mult_242_n21, mult_242_n20, mult_242_n19, 
      mult_242_n18, mult_242_n17, mult_242_n16, mult_242_n15, mult_242_n14, 
      mult_242_n13, mult_242_n12, mult_242_n11, mult_242_n10, mult_242_n9, 
      mult_242_n8, mult_242_n7, mult_242_n6, mult_242_n5, mult_242_n4, 
      mult_242_n3, mult_242_n2, mult_240_n130, mult_240_n129, mult_240_n128, 
      mult_240_n127, mult_240_n126, mult_240_n125, mult_240_n124, mult_240_n123
      , mult_240_n122, mult_240_n121, mult_240_n120, mult_240_n119, 
      mult_240_n70, mult_240_n69, mult_240_n68, mult_240_n67, mult_240_n65, 
      mult_240_n64, mult_240_n63, mult_240_n62, mult_240_n61, mult_240_n59, 
      mult_240_n58, mult_240_n57, mult_240_n56, mult_240_n55, mult_240_n54, 
      mult_240_n53, mult_240_n52, mult_240_n51, mult_240_n50, mult_240_n49, 
      mult_240_n48, mult_240_n47, mult_240_n46, mult_240_n44, mult_240_n43, 
      mult_240_n42, mult_240_n41, mult_240_n40, mult_240_n39, mult_240_n38, 
      mult_240_n37, mult_240_n36, mult_240_n35, mult_240_n34, mult_240_n32, 
      mult_240_n31, mult_240_n30, mult_240_n29, mult_240_n28, mult_240_n26, 
      mult_240_n25, mult_240_n24, mult_240_n23, mult_240_n22, mult_240_n21, 
      mult_240_n20, mult_240_n19, mult_240_n18, mult_240_n17, mult_240_n15, 
      mult_240_n14, mult_240_n12, mult_240_n11, mult_240_n10, mult_240_n9, 
      mult_240_n8, mult_240_n7, mult_240_n6, mult_240_n5, mult_240_n4, 
      mult_240_n3, mult_240_n2, mult_241_n179, mult_241_n178, mult_241_n177, 
      mult_241_n176, mult_241_n175, mult_241_n174, mult_241_n173, mult_241_n172
      , mult_241_n171, mult_241_n170, mult_241_n169, mult_241_n168, 
      mult_241_n167, mult_241_n115, mult_241_n114, mult_241_n113, mult_241_n112
      , mult_241_n111, mult_241_n110, mult_241_n109, mult_241_n108, 
      mult_241_n107, mult_241_n106, mult_241_n105, mult_241_n104, mult_241_n103
      , mult_241_n102, mult_241_n101, mult_241_n100, mult_241_n99, mult_241_n98
      , mult_241_n97, mult_241_n96, mult_241_n95, mult_241_n93, mult_241_n92, 
      mult_241_n91, mult_241_n90, mult_241_n89, mult_241_n88, mult_241_n87, 
      mult_241_n86, mult_241_n85, mult_241_n84, mult_241_n83, mult_241_n81, 
      mult_241_n80, mult_241_n79, mult_241_n78, mult_241_n77, mult_241_n76, 
      mult_241_n75, mult_241_n74, mult_241_n73, mult_241_n72, mult_241_n70, 
      mult_241_n69, mult_241_n68, mult_241_n67, mult_241_n66, mult_241_n65, 
      mult_241_n64, mult_241_n63, mult_241_n62, mult_241_n61, mult_241_n60, 
      mult_241_n59, mult_241_n58, mult_241_n57, mult_241_n56, mult_241_n55, 
      mult_241_n54, mult_241_n53, mult_241_n52, mult_241_n51, mult_241_n50, 
      mult_241_n49, mult_241_n48, mult_241_n47, mult_241_n46, mult_241_n45, 
      mult_241_n44, mult_241_n43, mult_241_n42, mult_241_n41, mult_241_n40, 
      mult_241_n39, mult_241_n38, mult_241_n37, mult_241_n36, mult_241_n35, 
      mult_241_n34, mult_241_n33, mult_241_n32, mult_241_n31, mult_241_n30, 
      mult_241_n29, mult_241_n28, mult_241_n27, mult_241_n26, mult_241_n25, 
      mult_241_n24, mult_241_n22, mult_241_n21, mult_241_n20, mult_241_n18, 
      mult_241_n17, mult_241_n16, mult_241_n15, mult_241_n14, mult_241_n13, 
      mult_241_n12, mult_241_n11, mult_241_n10, mult_241_n9, mult_241_n8, 
      mult_241_n7, mult_241_n6, mult_241_n5, mult_241_n4, mult_241_n3, 
      mult_241_n2, mult_239_n109, mult_239_n108, mult_239_n107, mult_239_n106, 
      mult_239_n105, mult_239_n104, mult_239_n103, mult_239_n102, mult_239_n101
      , mult_239_n100, mult_239_n99, mult_239_n98, mult_239_n96, mult_239_n47, 
      mult_239_n46, mult_239_n45, mult_239_n44, mult_239_n43, mult_239_n42, 
      mult_239_n41, mult_239_n40, mult_239_n39, mult_239_n38, mult_239_n37, 
      mult_239_n36, mult_239_n35, mult_239_n34, mult_239_n33, mult_239_n32, 
      mult_239_n31, mult_239_n30, mult_239_n29, mult_239_n28, mult_239_n27, 
      mult_239_n25, mult_239_n24, mult_239_n23, mult_239_n22, mult_239_n21, 
      mult_239_n19, mult_239_n17, mult_239_n15, mult_239_n13, mult_239_n12, 
      mult_239_n11, mult_239_n10, mult_239_n9, mult_239_n8, mult_239_n7, 
      mult_239_n6, mult_239_n5, mult_239_n4, mult_239_n3, mult_239_n2, 
      mult_239_n1 : std_logic;

begin
   
   U149 : OAI21D1 port map( A1 => n193, A2 => n247, B => n92, Z => n132);
   U150 : AOI22D1 port map( A1 => n190, A2 => a1_out_7_port, B1 => 
                           m2_out_14_port, B2 => n177, Z => n92);
   U151 : OAI21D1 port map( A1 => n193, A2 => n246, B => n94, Z => n133);
   U152 : AOI22D1 port map( A1 => n190, A2 => a1_out_6_port, B1 => 
                           m2_out_13_port, B2 => n177, Z => n94);
   U153 : OAI21D1 port map( A1 => n193, A2 => n245, B => n95, Z => n134);
   U154 : AOI22D1 port map( A1 => n190, A2 => a1_out_5_port, B1 => 
                           m2_out_12_port, B2 => n177, Z => n95);
   U155 : OAI21D1 port map( A1 => n193, A2 => n244, B => n96, Z => n135);
   U156 : AOI22D1 port map( A1 => n190, A2 => a1_out_4_port, B1 => 
                           m2_out_11_port, B2 => n177, Z => n96);
   U157 : OAI21D1 port map( A1 => n193, A2 => n243, B => n97, Z => n136);
   U158 : AOI22D1 port map( A1 => n190, A2 => a1_out_3_port, B1 => 
                           m2_out_10_port, B2 => n177, Z => n97);
   U159 : OAI21D1 port map( A1 => n193, A2 => n242, B => n98, Z => n137);
   U160 : AOI22D1 port map( A1 => n189, A2 => a1_out_2_port, B1 => 
                           m2_out_9_port, B2 => n177, Z => n98);
   U161 : OAI21D1 port map( A1 => n193, A2 => n241, B => n99, Z => n138);
   U162 : AOI22D1 port map( A1 => n189, A2 => a1_out_1_port, B1 => 
                           m2_out_8_port, B2 => n177, Z => n99);
   U163 : OAI21D1 port map( A1 => n193, A2 => n240, B => n100, Z => n139);
   U164 : AOI22D1 port map( A1 => n189, A2 => a1_out_0_port, B1 => 
                           m2_out_7_port, B2 => n177, Z => n100);
   U165 : OAI21D1 port map( A1 => n193, A2 => n239, B => n102, Z => n147);
   U166 : AOI22D1 port map( A1 => a2_out_7_port, A2 => n189, B1 => 
                           m4_out_14_port, B2 => n177, Z => n102);
   U167 : OAI21D1 port map( A1 => n193, A2 => n238, B => n103, Z => n148);
   U168 : AOI22D1 port map( A1 => a2_out_6_port, A2 => n189, B1 => 
                           m4_out_13_port, B2 => n177, Z => n103);
   U169 : OAI21D1 port map( A1 => n193, A2 => n237, B => n104, Z => n149);
   U170 : AOI22D1 port map( A1 => a2_out_5_port, A2 => n189, B1 => 
                           m4_out_12_port, B2 => n177, Z => n104);
   U171 : OAI21D1 port map( A1 => n193, A2 => n236, B => n105, Z => n150);
   U172 : AOI22D1 port map( A1 => a2_out_4_port, A2 => n189, B1 => 
                           m4_out_11_port, B2 => n177, Z => n105);
   U173 : OAI21D1 port map( A1 => n193, A2 => n235, B => n1060, Z => n151);
   U174 : AOI22D1 port map( A1 => a2_out_3_port, A2 => n189, B1 => 
                           m4_out_10_port, B2 => n177, Z => n1060);
   U175 : OAI21D1 port map( A1 => n193, A2 => n234, B => n1070, Z => n152);
   U176 : AOI22D1 port map( A1 => a2_out_2_port, A2 => n189, B1 => 
                           m4_out_9_port, B2 => n177, Z => n1070);
   U177 : OAI21D1 port map( A1 => n193, A2 => n233, B => n1080, Z => n153);
   U178 : AOI22D1 port map( A1 => a2_out_1_port, A2 => n189, B1 => 
                           m4_out_8_port, B2 => n177, Z => n1080);
   U179 : OAI21D1 port map( A1 => n193, A2 => n232, B => n1090, Z => n154);
   U180 : AOI22D1 port map( A1 => a2_out_0_port, A2 => n189, B1 => 
                           m4_out_7_port, B2 => n177, Z => n1090);
   U181 : OAI21D1 port map( A1 => n193, A2 => n217, B => n1120, Z => n162);
   U182 : AOI22D1 port map( A1 => m1_out_0_port, A2 => n189, B1 => 
                           m5_out_0_port, B2 => n177, Z => n1120);
   U183 : OAI21D1 port map( A1 => n193, A2 => n216, B => n1130, Z => n163);
   U184 : AOI22D1 port map( A1 => m1_out_1_port, A2 => n189, B1 => 
                           m5_out_1_port, B2 => n177, Z => n1130);
   U185 : OAI21D1 port map( A1 => n193, A2 => n215, B => n1140, Z => n164);
   U186 : AOI22D1 port map( A1 => m1_out_2_port, A2 => n189, B1 => 
                           m5_out_2_port, B2 => n177, Z => n1140);
   U187 : OAI21D1 port map( A1 => n193, A2 => n214, B => n1150, Z => n165);
   U188 : AOI22D1 port map( A1 => m1_out_3_port, A2 => n189, B1 => 
                           m5_out_3_port, B2 => n177, Z => n1150);
   U189 : OAI21D1 port map( A1 => n193, A2 => n213, B => n1160, Z => n166);
   U190 : AOI22D1 port map( A1 => m1_out_4_port, A2 => n189, B1 => 
                           m5_out_4_port, B2 => n177, Z => n1160);
   U191 : OAI21D1 port map( A1 => n193, A2 => n212, B => n1170, Z => n167);
   U192 : AOI22D1 port map( A1 => m1_out_5_port, A2 => n189, B1 => 
                           m5_out_5_port, B2 => n177, Z => n1170);
   U193 : OAI21D1 port map( A1 => n193, A2 => n211, B => n1180, Z => n168);
   U194 : AOI22D1 port map( A1 => m1_out_6_port, A2 => n189, B1 => 
                           m5_out_6_port, B2 => n177, Z => n1180);
   U195 : OAI21D1 port map( A1 => n193, A2 => n210, B => n1190, Z => n169);
   U196 : AOI22D1 port map( A1 => m1_out_7_port, A2 => n189, B1 => 
                           m5_out_7_port, B2 => n177, Z => n1190);
   U197 : OAI21D1 port map( A1 => n193, A2 => n209, B => n1200, Z => n170);
   U198 : AOI22D1 port map( A1 => m1_out_8_port, A2 => n189, B1 => 
                           m5_out_8_port, B2 => n177, Z => n1200);
   U199 : OAI21D1 port map( A1 => n193, A2 => n208, B => n1210, Z => n171);
   U200 : AOI22D1 port map( A1 => m1_out_9_port, A2 => n189, B1 => 
                           m5_out_9_port, B2 => n177, Z => n1210);
   U201 : OAI21D1 port map( A1 => n193, A2 => n207, B => n1220, Z => n172);
   U202 : AOI22D1 port map( A1 => m1_out_10_port, A2 => n189, B1 => 
                           m5_out_10_port, B2 => n177, Z => n1220);
   U203 : OAI21D1 port map( A1 => n193, A2 => n206, B => n1230, Z => n173);
   U204 : AOI22D1 port map( A1 => m1_out_11_port, A2 => n189, B1 => 
                           m5_out_11_port, B2 => n177, Z => n1230);
   U205 : OAI21D1 port map( A1 => n193, A2 => n205, B => n124, Z => n174);
   U206 : AOI22D1 port map( A1 => m1_out_12_port, A2 => n190, B1 => 
                           m5_out_12_port, B2 => n177, Z => n124);
   U207 : OAI21D1 port map( A1 => n193, A2 => n204, B => n125, Z => n175);
   U208 : AOI22D1 port map( A1 => m1_out_15, A2 => n189, B1 => m5_out_15, B2 =>
                           n177, Z => n125);
   U209 : OAI21D1 port map( A1 => n193, A2 => n203, B => n126, Z => n176);
   U210 : AOI22D1 port map( A1 => m1_out_15, A2 => n189, B1 => m5_out_15, B2 =>
                           n177, Z => n126);
   U211 : OAI22M10D1 port map( A1 => arx_r4_reg_9_port, A2 => n1110, B1 => n234
                           , B2 => n179, Z => a2_in_r_9_port);
   U212 : OAI22M10D1 port map( A1 => arx_r4_reg_8_port, A2 => n188, B1 => n233,
                           B2 => n179, Z => a2_in_r_8_port);
   U213 : OAI22M10D1 port map( A1 => arx_r4_reg_7_port, A2 => n188, B1 => n232,
                           B2 => n179, Z => a2_in_r_7_port);
   U214 : OAI22M10D1 port map( A1 => arx_r4_reg_6_port, A2 => n188, B1 => n225,
                           B2 => n179, Z => a2_in_r_6_port);
   U215 : OAI22M10D1 port map( A1 => arx_r4_reg_5_port, A2 => n188, B1 => n226,
                           B2 => n179, Z => a2_in_r_5_port);
   U216 : OAI22M10D1 port map( A1 => arx_r4_reg_4_port, A2 => n188, B1 => n227,
                           B2 => n179, Z => a2_in_r_4_port);
   U217 : OAI22M10D1 port map( A1 => arx_r4_reg_3_port, A2 => n188, B1 => n228,
                           B2 => n179, Z => a2_in_r_3_port);
   U218 : OAI22M10D1 port map( A1 => arx_r4_reg_2_port, A2 => n188, B1 => n229,
                           B2 => n179, Z => a2_in_r_2_port);
   U219 : OAI22M10D1 port map( A1 => arx_r4_reg_1_port, A2 => n188, B1 => n230,
                           B2 => n179, Z => a2_in_r_1_port);
   U220 : OAI22M10D1 port map( A1 => arx_r4_reg_14_port, A2 => n188, B1 => n239
                           , B2 => n179, Z => a2_in_r_14_port);
   U221 : OAI22M10D1 port map( A1 => arx_r4_reg_13_port, A2 => n1110, B1 => 
                           n238, B2 => n179, Z => a2_in_r_13_port);
   U222 : OAI22M10D1 port map( A1 => arx_r4_reg_12_port, A2 => n1110, B1 => 
                           n237, B2 => n179, Z => a2_in_r_12_port);
   U223 : OAI22M10D1 port map( A1 => arx_r4_reg_11_port, A2 => n1110, B1 => 
                           n236, B2 => n179, Z => a2_in_r_11_port);
   U224 : OAI22M10D1 port map( A1 => arx_r4_reg_10_port, A2 => n1110, B1 => 
                           n235, B2 => n179, Z => a2_in_r_10_port);
   U226 : OAI22D1 port map( A1 => n188, A2 => n234, B1 => n242, B2 => n179, Z 
                           => a1_in_r_9_port);
   U227 : OAI22D1 port map( A1 => n188, A2 => n233, B1 => n241, B2 => n179, Z 
                           => a1_in_r_8_port);
   U228 : OAI22D1 port map( A1 => n188, A2 => n232, B1 => n240, B2 => n179, Z 
                           => a1_in_r_7_port);
   U229 : OAI22D1 port map( A1 => n188, A2 => n225, B1 => n218, B2 => n179, Z 
                           => a1_in_r_6_port);
   U230 : OAI22D1 port map( A1 => n188, A2 => n226, B1 => n219, B2 => n179, Z 
                           => a1_in_r_5_port);
   U231 : OAI22D1 port map( A1 => n188, A2 => n227, B1 => n220, B2 => n179, Z 
                           => a1_in_r_4_port);
   U232 : OAI22D1 port map( A1 => n188, A2 => n228, B1 => n221, B2 => n179, Z 
                           => a1_in_r_3_port);
   U233 : OAI22D1 port map( A1 => n188, A2 => n229, B1 => n222, B2 => n179, Z 
                           => a1_in_r_2_port);
   U234 : OAI22D1 port map( A1 => n188, A2 => n230, B1 => n223, B2 => n179, Z 
                           => a1_in_r_1_port);
   U235 : OAI22D1 port map( A1 => n1110, A2 => n239, B1 => n247, B2 => n179, Z 
                           => a1_in_r_14_port);
   U236 : OAI22D1 port map( A1 => n1110, A2 => n238, B1 => n246, B2 => n179, Z 
                           => a1_in_r_13_port);
   U237 : OAI22D1 port map( A1 => n1110, A2 => n237, B1 => n245, B2 => n179, Z 
                           => a1_in_r_12_port);
   U238 : OAI22D1 port map( A1 => n1110, A2 => n236, B1 => n244, B2 => n179, Z 
                           => a1_in_r_11_port);
   U239 : OAI22D1 port map( A1 => n1110, A2 => n235, B1 => n243, B2 => n179, Z 
                           => a1_in_r_10_port);
   U240 : OAI22D1 port map( A1 => n188, A2 => n231, B1 => n224, B2 => n179, Z 
                           => a1_in_r_0_port);
   U241 : OAI22M10D1 port map( A1 => arx_i1_reg_2_port, A2 => n179, B1 => n1110
                           , B2 => n242, Z => a1_in_l_9_port);
   U242 : OAI22M10D1 port map( A1 => arx_i1_reg_1_port, A2 => n179, B1 => n1110
                           , B2 => n241, Z => a1_in_l_8_port);
   U243 : OAI22M10D1 port map( A1 => arx_i1_reg_0_port, A2 => n179, B1 => n188,
                           B2 => n240, Z => a1_in_l_7_port);
   U244 : OAI22M10D1 port map( A1 => arx_i1_reg_7_port, A2 => n179, B1 => n1110
                           , B2 => n247, Z => a1_in_l_14_port);
   U245 : OAI22M10D1 port map( A1 => arx_i1_reg_6_port, A2 => n179, B1 => n1110
                           , B2 => n246, Z => a1_in_l_13_port);
   U246 : OAI22M10D1 port map( A1 => arx_i1_reg_5_port, A2 => n179, B1 => n1110
                           , B2 => n245, Z => a1_in_l_12_port);
   U247 : OAI22M10D1 port map( A1 => arx_i1_reg_4_port, A2 => n179, B1 => n1110
                           , B2 => n244, Z => a1_in_l_11_port);
   U248 : OAI22M10D1 port map( A1 => arx_i1_reg_3_port, A2 => n179, B1 => n1110
                           , B2 => n243, Z => a1_in_l_10_port);
   arx_r1_reg_reg_14 : DFFRPQ1 port map( D => n176, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_14_port);
   arx_r4_reg_reg_14 : DFERPQ1 port map( D => m3_out_14_port, CEB => n1100, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_14_port);
   arx_i1_reg_reg_7 : DFERPQ1 port map( D => data_in(7), CEB => n127, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_7_port);
   arx_r2_reg_reg_14 : DFFRPQ1 port map( D => n132, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_14_port);
   arx_r3_reg_reg_14 : DFFRPQ1 port map( D => n147, CK => clock, RB => resetn, 
                           Q => arx_r3_reg_14_port);
   arx_r1_reg_reg_13 : DFFRPQ1 port map( D => n175, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_13_port);
   arx_r4_reg_reg_13 : DFERPQ1 port map( D => m3_out_13_port, CEB => n1100, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_13_port);
   arx_i1_reg_reg_6 : DFERPQ1 port map( D => data_in(6), CEB => n127, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_6_port);
   arx_r2_reg_reg_13 : DFFRPQ1 port map( D => n133, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_13_port);
   arx_r3_reg_reg_13 : DFFRPQ1 port map( D => n148, CK => clock, RB => resetn, 
                           Q => arx_r3_reg_13_port);
   arx_r1_reg_reg_12 : DFFRPQ1 port map( D => n174, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_12_port);
   arx_r4_reg_reg_12 : DFERPQ1 port map( D => m3_out_12_port, CEB => n1100, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_12_port);
   arx_i1_reg_reg_5 : DFERPQ1 port map( D => data_in(5), CEB => n127, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_5_port);
   arx_r2_reg_reg_12 : DFFRPQ1 port map( D => n134, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_12_port);
   arx_r3_reg_reg_12 : DFFRPQ1 port map( D => n149, CK => clock, RB => resetn, 
                           Q => arx_r3_reg_12_port);
   arx_r1_reg_reg_11 : DFFRPQ1 port map( D => n173, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_11_port);
   arx_r4_reg_reg_11 : DFERPQ1 port map( D => m3_out_11_port, CEB => n1100, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_11_port);
   arx_i1_reg_reg_4 : DFERPQ1 port map( D => data_in(4), CEB => n127, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_4_port);
   arx_r2_reg_reg_11 : DFFRPQ1 port map( D => n135, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_11_port);
   arx_r3_reg_reg_11 : DFFRPQ1 port map( D => n150, CK => clock, RB => resetn, 
                           Q => arx_r3_reg_11_port);
   arx_r1_reg_reg_10 : DFFRPQ1 port map( D => n172, CK => clock, RB => resetn, 
                           Q => arx_r1_reg_10_port);
   arx_r4_reg_reg_10 : DFERPQ1 port map( D => m3_out_10_port, CEB => n1100, CK 
                           => clock, RB => resetn, Q => arx_r4_reg_10_port);
   arx_i1_reg_reg_3 : DFERPQ1 port map( D => data_in(3), CEB => n127, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_3_port);
   arx_r2_reg_reg_10 : DFFRPQ1 port map( D => n136, CK => clock, RB => resetn, 
                           Q => arx_r2_reg_10_port);
   arx_r3_reg_reg_10 : DFFRPQ1 port map( D => n151, CK => clock, RB => resetn, 
                           Q => arx_r3_reg_10_port);
   arx_r1_reg_reg_9 : DFFRPQ1 port map( D => n171, CK => clock, RB => resetn, Q
                           => arx_r1_reg_9_port);
   arx_r4_reg_reg_9 : DFERPQ1 port map( D => m3_out_9_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_9_port);
   arx_i1_reg_reg_2 : DFERPQ1 port map( D => data_in(2), CEB => n127, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_2_port);
   arx_r2_reg_reg_9 : DFFRPQ1 port map( D => n137, CK => clock, RB => resetn, Q
                           => arx_r2_reg_9_port);
   arx_r3_reg_reg_9 : DFFRPQ1 port map( D => n152, CK => clock, RB => resetn, Q
                           => arx_r3_reg_9_port);
   arx_r1_reg_reg_8 : DFFRPQ1 port map( D => n170, CK => clock, RB => resetn, Q
                           => arx_r1_reg_8_port);
   arx_r4_reg_reg_8 : DFERPQ1 port map( D => m3_out_8_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_8_port);
   arx_i1_reg_reg_1 : DFERPQ1 port map( D => data_in(1), CEB => n127, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_1_port);
   arx_r2_reg_reg_8 : DFFRPQ1 port map( D => n138, CK => clock, RB => resetn, Q
                           => arx_r2_reg_8_port);
   arx_r3_reg_reg_8 : DFFRPQ1 port map( D => n153, CK => clock, RB => resetn, Q
                           => arx_r3_reg_8_port);
   arx_r1_reg_reg_7 : DFFRPQ1 port map( D => n169, CK => clock, RB => resetn, Q
                           => arx_r1_reg_7_port);
   arx_r4_reg_reg_7 : DFERPQ1 port map( D => m3_out_7_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_7_port);
   arx_i1_reg_reg_0 : DFERPQ1 port map( D => data_in(0), CEB => n127, CK => 
                           clock, RB => resetn, Q => arx_i1_reg_0_port);
   arx_r2_reg_reg_7 : DFFRPQ1 port map( D => n139, CK => clock, RB => resetn, Q
                           => arx_r2_reg_7_port);
   arx_r3_reg_reg_7 : DFFRPQ1 port map( D => n154, CK => clock, RB => resetn, Q
                           => arx_r3_reg_7_port);
   arx_d1_reg_reg_14 : DFERPQ1 port map( D => a1_out_7_port, CEB => n178, CK =>
                           clock, RB => resetn, Q => arx_d1_reg_14_port);
   arx_d3_reg_reg_14 : DFERPQ1 port map( D => arx_d2_reg_14_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => N51);
   arx_d3_reg_reg_13 : DFERPQ1 port map( D => arx_d2_reg_13_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => N50);
   arx_d1_reg_reg_13 : DFERPQ1 port map( D => a1_out_6_port, CEB => n178, CK =>
                           clock, RB => resetn, Q => arx_d1_reg_13_port);
   arx_r1_reg_reg_6 : DFFRPQ1 port map( D => n168, CK => clock, RB => resetn, Q
                           => arx_r1_reg_6_port);
   arx_r4_reg_reg_6 : DFERPQ1 port map( D => m3_out_6_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_6_port);
   arx_r2_reg_reg_6 : DFFRPQ1 port map( D => n140, CK => clock, RB => resetn, Q
                           => arx_r2_reg_6_port);
   arx_d1_reg_reg_12 : DFERPQ1 port map( D => a1_out_5_port, CEB => n178, CK =>
                           clock, RB => resetn, Q => arx_d1_reg_12_port);
   arx_r3_reg_reg_6 : DFFRPQ1 port map( D => n155, CK => clock, RB => resetn, Q
                           => arx_r3_reg_6_port);
   arx_r4_reg_reg_5 : DFERPQ1 port map( D => m3_out_5_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_5_port);
   arx_r1_reg_reg_5 : DFFRPQ1 port map( D => n167, CK => clock, RB => resetn, Q
                           => arx_r1_reg_5_port);
   arx_d3_reg_reg_12 : DFERPQ1 port map( D => arx_d2_reg_12_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => N49);
   arx_r2_reg_reg_5 : DFFRPQ1 port map( D => n141, CK => clock, RB => resetn, Q
                           => arx_r2_reg_5_port);
   arx_r3_reg_reg_5 : DFFRPQ1 port map( D => n156, CK => clock, RB => resetn, Q
                           => arx_r3_reg_5_port);
   arx_d3_reg_reg_9 : DFERPQ1 port map( D => arx_d2_reg_9_port, CEB => n178, CK
                           => clock, RB => resetn, Q => N46);
   arx_d1_reg_reg_11 : DFERPQ1 port map( D => a1_out_4_port, CEB => n178, CK =>
                           clock, RB => resetn, Q => arx_d1_reg_11_port);
   arx_d3_reg_reg_8 : DFERPQ1 port map( D => arx_d2_reg_8_port, CEB => n178, CK
                           => clock, RB => resetn, Q => N45);
   arx_d3_reg_reg_10 : DFERPQ1 port map( D => arx_d2_reg_10_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => N47);
   arx_d3_reg_reg_11 : DFERPQ1 port map( D => arx_d2_reg_11_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => N48);
   arx_d3_reg_reg_7 : DFERPQ1 port map( D => arx_d2_reg_7_port, CEB => n178, CK
                           => clock, RB => resetn, Q => N44);
   arx_r4_reg_reg_4 : DFERPQ1 port map( D => m3_out_4_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_4_port);
   arx_r1_reg_reg_4 : DFFRPQ1 port map( D => n166, CK => clock, RB => resetn, Q
                           => arx_r1_reg_4_port);
   arx_d1_reg_reg_10 : DFERPQ1 port map( D => a1_out_3_port, CEB => n178, CK =>
                           clock, RB => resetn, Q => arx_d1_reg_10_port);
   arx_r2_reg_reg_4 : DFFRPQ1 port map( D => n142, CK => clock, RB => resetn, Q
                           => arx_r2_reg_4_port);
   arx_r3_reg_reg_4 : DFFRPQ1 port map( D => n157, CK => clock, RB => resetn, Q
                           => arx_r3_reg_4_port);
   arx_r4_reg_reg_3 : DFERPQ1 port map( D => m3_out_3_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_3_port);
   arx_r1_reg_reg_3 : DFFRPQ1 port map( D => n165, CK => clock, RB => resetn, Q
                           => arx_r1_reg_3_port);
   arx_r2_reg_reg_3 : DFFRPQ1 port map( D => n143, CK => clock, RB => resetn, Q
                           => arx_r2_reg_3_port);
   arx_r3_reg_reg_3 : DFFRPQ1 port map( D => n158, CK => clock, RB => resetn, Q
                           => arx_r3_reg_3_port);
   arx_d2_reg_reg_14 : DFERPQ1 port map( D => arx_d1_reg_14_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d2_reg_14_port);
   arx_d1_reg_reg_9 : DFERPQ1 port map( D => a1_out_2_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => arx_d1_reg_9_port);
   arx_d1_reg_reg_8 : DFERPQ1 port map( D => a1_out_1_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => arx_d1_reg_8_port);
   arx_d1_reg_reg_7 : DFERPQ1 port map( D => a1_out_0_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => arx_d1_reg_7_port);
   arx_r4_reg_reg_2 : DFERPQ1 port map( D => m3_out_2_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_2_port);
   arx_r1_reg_reg_2 : DFFRPQ1 port map( D => n164, CK => clock, RB => resetn, Q
                           => arx_r1_reg_2_port);
   arx_r2_reg_reg_2 : DFFRPQ1 port map( D => n144, CK => clock, RB => resetn, Q
                           => arx_r2_reg_2_port);
   arx_r3_reg_reg_2 : DFFRPQ1 port map( D => n159, CK => clock, RB => resetn, Q
                           => arx_r3_reg_2_port);
   arx_d2_reg_reg_12 : DFERPQ1 port map( D => arx_d1_reg_12_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d2_reg_12_port);
   arx_d2_reg_reg_13 : DFERPQ1 port map( D => arx_d1_reg_13_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d2_reg_13_port);
   arx_r1_reg_reg_0 : DFFRPQ1 port map( D => n162, CK => clock, RB => resetn, Q
                           => arx_r1_reg_0_port);
   arx_r2_reg_reg_0 : DFFRPQ1 port map( D => n146, CK => clock, RB => resetn, Q
                           => arx_r2_reg_0_port);
   arx_r1_reg_reg_1 : DFFRPQ1 port map( D => n163, CK => clock, RB => resetn, Q
                           => arx_r1_reg_1_port);
   arx_r3_reg_reg_0 : DFFRPQ1 port map( D => n161, CK => clock, RB => resetn, Q
                           => arx_r3_reg_0_port);
   arx_r4_reg_reg_1 : DFERPQ1 port map( D => m3_out_1_port, CEB => n1100, CK =>
                           clock, RB => resetn, Q => arx_r4_reg_1_port);
   arx_d2_reg_reg_11 : DFERPQ1 port map( D => arx_d1_reg_11_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d2_reg_11_port);
   arx_r2_reg_reg_1 : DFFRPQ1 port map( D => n145, CK => clock, RB => resetn, Q
                           => arx_r2_reg_1_port);
   arx_r3_reg_reg_1 : DFFRPQ1 port map( D => n160, CK => clock, RB => resetn, Q
                           => arx_r3_reg_1_port);
   arx_d2_reg_reg_10 : DFERPQ1 port map( D => arx_d1_reg_10_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d2_reg_10_port);
   arx_d2_reg_reg_7 : DFERPQ1 port map( D => arx_d1_reg_7_port, CEB => n178, CK
                           => clock, RB => resetn, Q => arx_d2_reg_7_port);
   arx_d2_reg_reg_8 : DFERPQ1 port map( D => arx_d1_reg_8_port, CEB => n178, CK
                           => clock, RB => resetn, Q => arx_d2_reg_8_port);
   arx_d2_reg_reg_9 : DFERPQ1 port map( D => arx_d1_reg_9_port, CEB => n178, CK
                           => clock, RB => resetn, Q => arx_d2_reg_9_port);
   arx_state_reg_reg_1 : DFFRPQ1 port map( D => n193, CK => clock, RB => resetn
                           , Q => arx_state_reg_1_port);
   arx_state_reg_reg_0 : DFFRPQ1 port map( D => state_0, CK => clock, RB => 
                           resetn, Q => arx_state_reg_0_port);
   arx_o1_reg_reg_7 : DFERPQ1 port map( D => a2_out_7_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => data_out(7));
   arx_o1_reg_reg_0 : DFERPQ1 port map( D => a2_out_0_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => data_out(0));
   arx_o1_reg_reg_1 : DFERPQ1 port map( D => a2_out_1_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => data_out(1));
   arx_o1_reg_reg_2 : DFERPQ1 port map( D => a2_out_2_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => data_out(2));
   arx_o1_reg_reg_3 : DFERPQ1 port map( D => a2_out_3_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => data_out(3));
   arx_o1_reg_reg_4 : DFERPQ1 port map( D => a2_out_4_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => data_out(4));
   arx_o1_reg_reg_5 : DFERPQ1 port map( D => a2_out_5_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => data_out(5));
   arx_o1_reg_reg_6 : DFERPQ1 port map( D => a2_out_6_port, CEB => n178, CK => 
                           clock, RB => resetn, Q => data_out(6));
   U249 : INVBD2 port map( A => arx_d2_reg_14_port, Z => n187);
   U250 : INVBD2 port map( A => arx_d2_reg_13_port, Z => n185);
   U251 : INVBD2 port map( A => arx_d2_reg_12_port, Z => n186);
   U252 : INVBD2 port map( A => arx_d2_reg_11_port, Z => n184);
   U253 : INVBD2 port map( A => arx_d2_reg_10_port, Z => n182);
   U254 : INVBD2 port map( A => arx_d2_reg_9_port, Z => n180);
   U255 : INVBD2 port map( A => arx_d2_reg_8_port, Z => n181);
   U256 : INVBD2 port map( A => arx_d2_reg_7_port, Z => n183);
   U257 : NOR2D2 port map( A1 => n231, A2 => n179, Z => a2_in_r_0_port);
   U258 : NOR2D2 port map( A1 => n202, A2 => arx_state_reg_1_port, Z => n177);
   U259 : OR2D1 port map( A1 => n177, A2 => state_0, Z => n178);
   U260 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => 
                           arx_state_reg_1_port, Z => n179);
   U261 : INVD1 port map( A => n191, Z => n193);
   U262 : INVD1 port map( A => n192, Z => n191);
   U263 : INVD1 port map( A => n101, Z => n192);
   U264 : NAN2D1 port map( A1 => n193, A2 => n188, Z => n1100);
   U265 : INVD1 port map( A => m5_in_l_0, Z => n194);
   U266 : NOR2M1D1 port map( A1 => n179, A2 => n190, Z => n130);
   U267 : INVD1 port map( A => n189, Z => n188);
   U268 : NOR2D1 port map( A1 => n177, A2 => n190, Z => n101);
   U269 : NAN2D1 port map( A1 => n101, A2 => n179, Z => n127);
   U270 : NAN2M1D1 port map( A1 => n177, A2 => n129, Z => m5_in_l_0);
   U271 : NOR2D1 port map( A1 => n130, A2 => n216, Z => a2_in_l_1_port);
   U272 : NOR2D1 port map( A1 => n130, A2 => n217, Z => a2_in_l_0_port);
   U273 : INVD1 port map( A => n1110, Z => n190);
   U274 : NOR2D1 port map( A1 => n188, A2 => n224, Z => a1_in_l_0_port);
   U275 : NOR2D1 port map( A1 => n188, A2 => n218, Z => a1_in_l_6_port);
   U276 : NOR2D1 port map( A1 => n188, A2 => n222, Z => a1_in_l_2_port);
   U277 : NOR2D1 port map( A1 => n188, A2 => n221, Z => a1_in_l_3_port);
   U278 : NOR2D1 port map( A1 => n188, A2 => n220, Z => a1_in_l_4_port);
   U279 : INVD1 port map( A => n1110, Z => n189);
   U280 : NOR2D1 port map( A1 => n194, A2 => n248, Z => m2_in_r_0_port);
   U281 : NOR2D1 port map( A1 => n194, A2 => n201, Z => m2_in_r_1_port);
   U282 : NOR2D1 port map( A1 => n188, A2 => n223, Z => a1_in_l_1_port);
   U283 : NOR2D1 port map( A1 => n194, A2 => n200, Z => m2_in_r_2_port);
   U284 : NOR2D1 port map( A1 => n194, A2 => n199, Z => m2_in_r_3_port);
   U285 : NOR2D1 port map( A1 => n191, A2 => n198, Z => m1_in_r_4_port);
   U286 : NOR2D1 port map( A1 => n191, A2 => n199, Z => m1_in_r_3_port);
   U287 : NOR2D1 port map( A1 => n191, A2 => n248, Z => m1_in_r_0_port);
   U288 : NOR2D1 port map( A1 => n191, A2 => n201, Z => m1_in_r_1_port);
   U289 : NOR2D1 port map( A1 => n191, A2 => n200, Z => m1_in_r_2_port);
   U290 : NOR2D1 port map( A1 => n191, A2 => n197, Z => m1_in_r_5_port);
   U291 : NOR2D1 port map( A1 => n130, A2 => n212, Z => a2_in_l_5_port);
   U292 : NOR2D1 port map( A1 => n194, A2 => n198, Z => m2_in_r_4_port);
   U293 : NOR2D1 port map( A1 => n194, A2 => n196, Z => m2_in_r_6_port);
   U294 : NOR2D1 port map( A1 => n194, A2 => n197, Z => m2_in_r_5_port);
   U295 : NOR2D1 port map( A1 => n101, A2 => n196, Z => m1_in_r_6_port);
   U296 : NOR2D1 port map( A1 => n101, A2 => n195, Z => m1_in_r_7_port);
   U297 : NOR2D1 port map( A1 => n188, A2 => n219, Z => a1_in_l_5_port);
   U298 : NOR2D1 port map( A1 => n194, A2 => n195, Z => m2_in_r_7_port);
   U299 : NOR2D1 port map( A1 => n130, A2 => n203, Z => a2_in_l_14_port);
   U300 : NAN2D1 port map( A1 => n188, A2 => n129, Z => state_0);
   U301 : INVD1 port map( A => arx_state_reg_0_port, Z => n202);
   U302 : NOR2D1 port map( A1 => n180, A2 => n194, Z => m4_in_r_2_port);
   U303 : NOR2D1 port map( A1 => n181, A2 => n194, Z => m4_in_r_1_port);
   U304 : NOR2D1 port map( A1 => n182, A2 => n194, Z => m4_in_r_3_port);
   U305 : NOR2D1 port map( A1 => n183, A2 => n194, Z => m4_in_r_0_port);
   U306 : NAN2M1D1 port map( A1 => arx_state_reg_1_port, A2 => n202, Z => n129)
                           ;
   U307 : NOR2D1 port map( A1 => n130, A2 => n211, Z => a2_in_l_6_port);
   U308 : NOR2D1 port map( A1 => n130, A2 => n210, Z => a2_in_l_7_port);
   U309 : NOR2D1 port map( A1 => n130, A2 => n209, Z => a2_in_l_8_port);
   U310 : NOR2D1 port map( A1 => n130, A2 => n208, Z => a2_in_l_9_port);
   U311 : NOR2D1 port map( A1 => n130, A2 => n207, Z => a2_in_l_10_port);
   U312 : NOR2D1 port map( A1 => n130, A2 => n206, Z => a2_in_l_11_port);
   U313 : NOR2D1 port map( A1 => n130, A2 => n205, Z => a2_in_l_12_port);
   U314 : NOR2D1 port map( A1 => n130, A2 => n204, Z => a2_in_l_13_port);
   U315 : NOR2D1 port map( A1 => n130, A2 => n215, Z => a2_in_l_2_port);
   U316 : NOR2D1 port map( A1 => n130, A2 => n214, Z => a2_in_l_3_port);
   U317 : NOR2D1 port map( A1 => n130, A2 => n213, Z => a2_in_l_4_port);
   U318 : NOR2D1 port map( A1 => n184, A2 => n194, Z => m4_in_r_4_port);
   U319 : NAN2D1 port map( A1 => arx_state_reg_1_port, A2 => n202, Z => n1110);
   U320 : NOR2D1 port map( A1 => n185, A2 => n194, Z => m4_in_r_6_port);
   U321 : NOR2D1 port map( A1 => n186, A2 => n194, Z => m4_in_r_5_port);
   U322 : AND2D1 port map( A1 => N48, A2 => m5_in_l_0, Z => m5_in_r_4_port);
   U323 : AND2D1 port map( A1 => N45, A2 => m5_in_l_0, Z => m5_in_r_1_port);
   U324 : AND2D1 port map( A1 => N46, A2 => m5_in_l_0, Z => m5_in_r_2_port);
   U325 : AND2D1 port map( A1 => N47, A2 => m5_in_l_0, Z => m5_in_r_3_port);
   U326 : AND2D1 port map( A1 => N44, A2 => m5_in_l_0, Z => m5_in_r_0_port);
   U327 : NOR2D1 port map( A1 => n187, A2 => n194, Z => m4_in_r_7_port);
   U328 : AND2D1 port map( A1 => N49, A2 => m5_in_l_0, Z => m5_in_r_5_port);
   U329 : AND2D1 port map( A1 => N50, A2 => m5_in_l_0, Z => m5_in_r_6_port);
   U330 : AND2D1 port map( A1 => N51, A2 => m5_in_l_0, Z => m5_in_r_7_port);
   U331 : INVD1 port map( A => arx_r3_reg_1_port, Z => n230);
   U332 : INVD1 port map( A => arx_r2_reg_1_port, Z => n223);
   U333 : INVD1 port map( A => arx_r3_reg_0_port, Z => n231);
   U334 : INVD1 port map( A => arx_r1_reg_1_port, Z => n216);
   U335 : INVD1 port map( A => arx_r2_reg_0_port, Z => n224);
   U336 : INVD1 port map( A => arx_r1_reg_0_port, Z => n217);
   U337 : INVD1 port map( A => arx_r3_reg_2_port, Z => n229);
   U338 : INVD1 port map( A => arx_r2_reg_2_port, Z => n222);
   U339 : INVD1 port map( A => arx_r1_reg_2_port, Z => n215);
   U340 : INVD1 port map( A => arx_d1_reg_7_port, Z => n248);
   U341 : INVD1 port map( A => arx_d1_reg_8_port, Z => n201);
   U342 : INVD1 port map( A => arx_d1_reg_9_port, Z => n200);
   U343 : INVD1 port map( A => arx_r3_reg_3_port, Z => n228);
   U344 : AO22D1 port map( A1 => m4_out_6_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_6_port, Z => n155);
   U345 : INVD1 port map( A => arx_r2_reg_3_port, Z => n221);
   U346 : INVD1 port map( A => arx_r1_reg_3_port, Z => n214);
   U347 : AO22D1 port map( A1 => m2_out_6_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_6_port, Z => n140);
   U348 : INVD1 port map( A => arx_r3_reg_4_port, Z => n227);
   U349 : INVD1 port map( A => arx_r2_reg_4_port, Z => n220);
   U350 : INVD1 port map( A => arx_d1_reg_10_port, Z => n199);
   U351 : INVD1 port map( A => arx_r1_reg_4_port, Z => n213);
   U352 : AO22D1 port map( A1 => m4_out_5_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_5_port, Z => n156);
   U353 : INVD1 port map( A => arx_d1_reg_11_port, Z => n198);
   U354 : INVD1 port map( A => arx_r3_reg_5_port, Z => n226);
   U355 : INVD1 port map( A => arx_r2_reg_5_port, Z => n219);
   U356 : AO22D1 port map( A1 => m2_out_5_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_5_port, Z => n141);
   U357 : INVD1 port map( A => arx_r1_reg_5_port, Z => n212);
   U358 : INVD1 port map( A => arx_r3_reg_6_port, Z => n225);
   U359 : AO22D1 port map( A1 => m4_out_4_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_4_port, Z => n157);
   U360 : INVD1 port map( A => arx_d1_reg_12_port, Z => n197);
   U361 : INVD1 port map( A => arx_r2_reg_6_port, Z => n218);
   U362 : INVD1 port map( A => arx_r1_reg_6_port, Z => n211);
   U363 : INVD1 port map( A => arx_d1_reg_13_port, Z => n196);
   U364 : AO22D1 port map( A1 => m2_out_4_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_4_port, Z => n142);
   U365 : INVD1 port map( A => arx_d1_reg_14_port, Z => n195);
   U366 : AO22D1 port map( A1 => m4_out_3_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_3_port, Z => n158);
   U367 : INVD1 port map( A => arx_r3_reg_7_port, Z => n232);
   U368 : INVD1 port map( A => arx_r2_reg_7_port, Z => n240);
   U369 : INVD1 port map( A => arx_r1_reg_7_port, Z => n210);
   U370 : AO22D1 port map( A1 => m2_out_3_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_3_port, Z => n143);
   U371 : INVD1 port map( A => arx_r3_reg_8_port, Z => n233);
   U372 : INVD1 port map( A => arx_r2_reg_8_port, Z => n241);
   U373 : AO22D1 port map( A1 => m4_out_2_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_2_port, Z => n159);
   U374 : INVD1 port map( A => arx_r1_reg_8_port, Z => n209);
   U375 : AO22D1 port map( A1 => m2_out_2_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_2_port, Z => n144);
   U376 : INVD1 port map( A => arx_r3_reg_9_port, Z => n234);
   U377 : INVD1 port map( A => arx_r2_reg_9_port, Z => n242);
   U378 : INVD1 port map( A => arx_r1_reg_9_port, Z => n208);
   U379 : AO22D1 port map( A1 => m4_out_1_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_1_port, Z => n160);
   U380 : AO22D1 port map( A1 => m2_out_1_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_1_port, Z => n145);
   U381 : INVD1 port map( A => arx_r3_reg_10_port, Z => n235);
   U382 : INVD1 port map( A => arx_r2_reg_10_port, Z => n243);
   U383 : INVD1 port map( A => arx_r1_reg_10_port, Z => n207);
   U384 : AO22D1 port map( A1 => m2_out_0_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_0_port, Z => n146);
   U385 : AO22D1 port map( A1 => m4_out_0_port, A2 => n177, B1 => n191, B2 => 
                           arx_r3_reg_0_port, Z => n161);
   U386 : INVD1 port map( A => arx_r3_reg_11_port, Z => n236);
   U387 : INVD1 port map( A => arx_r2_reg_11_port, Z => n244);
   U388 : INVD1 port map( A => arx_r1_reg_11_port, Z => n206);
   U389 : INVD1 port map( A => arx_r3_reg_12_port, Z => n237);
   U390 : INVD1 port map( A => arx_r2_reg_12_port, Z => n245);
   U391 : INVD1 port map( A => arx_r1_reg_12_port, Z => n205);
   U392 : INVD1 port map( A => arx_r3_reg_13_port, Z => n238);
   U393 : INVD1 port map( A => arx_r2_reg_13_port, Z => n246);
   U394 : INVD1 port map( A => arx_r1_reg_13_port, Z => n204);
   U395 : INVD1 port map( A => arx_r3_reg_14_port, Z => n239);
   U396 : INVD1 port map( A => arx_r2_reg_14_port, Z => n247);
   U397 : INVD1 port map( A => arx_r1_reg_14_port, Z => n203);
   U398 : TIELO port map( Z => net1801);
   U399 : EXOR2D1 port map( A1 => N114, A2 => add_416_C243_rn_carry_7_port, Z 
                           => a1_out_7_port);
   U400 : AND2D1 port map( A1 => add_416_C243_rn_carry_6_port, A2 => N113, Z =>
                           add_416_C243_rn_carry_7_port);
   U401 : EXOR2D1 port map( A1 => N113, A2 => add_416_C243_rn_carry_6_port, Z 
                           => a1_out_6_port);
   U402 : AND2D1 port map( A1 => add_416_C243_rn_carry_5_port, A2 => N112, Z =>
                           add_416_C243_rn_carry_6_port);
   U403 : EXOR2D1 port map( A1 => N112, A2 => add_416_C243_rn_carry_5_port, Z 
                           => a1_out_5_port);
   U404 : AND2D1 port map( A1 => add_416_C243_rn_carry_4_port, A2 => N111, Z =>
                           add_416_C243_rn_carry_5_port);
   U405 : EXOR2D1 port map( A1 => N111, A2 => add_416_C243_rn_carry_4_port, Z 
                           => a1_out_4_port);
   U406 : AND2D1 port map( A1 => add_416_C243_rn_carry_3_port, A2 => N110, Z =>
                           add_416_C243_rn_carry_4_port);
   U407 : EXOR2D1 port map( A1 => N110, A2 => add_416_C243_rn_carry_3_port, Z 
                           => a1_out_3_port);
   U408 : AND2D1 port map( A1 => add_416_C243_rn_carry_2_port, A2 => N109, Z =>
                           add_416_C243_rn_carry_3_port);
   U409 : EXOR2D1 port map( A1 => N109, A2 => add_416_C243_rn_carry_2_port, Z 
                           => a1_out_2_port);
   U410 : AND2D1 port map( A1 => add_416_C243_rn_carry_1_port, A2 => N108, Z =>
                           add_416_C243_rn_carry_2_port);
   U411 : EXOR2D1 port map( A1 => N108, A2 => add_416_C243_rn_carry_1_port, Z 
                           => a1_out_1_port);
   U412 : AND2D1 port map( A1 => N107, A2 => N106, Z => 
                           add_416_C243_rn_carry_1_port);
   U413 : EXOR2D1 port map( A1 => N106, A2 => N107, Z => a1_out_0_port);
   U414 : EXOR2D1 port map( A1 => N123, A2 => add_416_C244_rn_carry_7_port, Z 
                           => a2_out_7_port);
   U415 : AND2D1 port map( A1 => add_416_C244_rn_carry_6_port, A2 => N122, Z =>
                           add_416_C244_rn_carry_7_port);
   U416 : EXOR2D1 port map( A1 => N122, A2 => add_416_C244_rn_carry_6_port, Z 
                           => a2_out_6_port);
   U417 : AND2D1 port map( A1 => add_416_C244_rn_carry_5_port, A2 => N121, Z =>
                           add_416_C244_rn_carry_6_port);
   U418 : EXOR2D1 port map( A1 => N121, A2 => add_416_C244_rn_carry_5_port, Z 
                           => a2_out_5_port);
   U419 : AND2D1 port map( A1 => add_416_C244_rn_carry_4_port, A2 => N120, Z =>
                           add_416_C244_rn_carry_5_port);
   U420 : EXOR2D1 port map( A1 => N120, A2 => add_416_C244_rn_carry_4_port, Z 
                           => a2_out_4_port);
   U421 : AND2D1 port map( A1 => add_416_C244_rn_carry_3_port, A2 => N119, Z =>
                           add_416_C244_rn_carry_4_port);
   U422 : EXOR2D1 port map( A1 => N119, A2 => add_416_C244_rn_carry_3_port, Z 
                           => a2_out_3_port);
   U423 : AND2D1 port map( A1 => add_416_C244_rn_carry_2_port, A2 => N118, Z =>
                           add_416_C244_rn_carry_3_port);
   U424 : EXOR2D1 port map( A1 => N118, A2 => add_416_C244_rn_carry_2_port, Z 
                           => a2_out_2_port);
   U425 : AND2D1 port map( A1 => add_416_C244_rn_carry_1_port, A2 => N117, Z =>
                           add_416_C244_rn_carry_2_port);
   U426 : EXOR2D1 port map( A1 => N117, A2 => add_416_C244_rn_carry_1_port, Z 
                           => a2_out_1_port);
   U427 : AND2D1 port map( A1 => N116, A2 => N115, Z => 
                           add_416_C244_rn_carry_1_port);
   U428 : EXOR2D1 port map( A1 => N115, A2 => N116, Z => a2_out_0_port);
   add_244_U10 : OAI211D1 port map( A1 => a2_in_l_1_port, A2 => a2_in_r_1_port,
                           B => a2_in_l_0_port, C => a2_in_r_0_port, Z => 
                           add_244_n9);
   add_244_U9 : OAI21M20D1 port map( A1 => a2_in_l_1_port, A2 => a2_in_r_1_port
                           , B => add_244_n9, Z => add_244_n7);
   add_244_U8 : OAI21D1 port map( A1 => a2_in_l_2_port, A2 => add_244_n7, B => 
                           a2_in_r_2_port, Z => add_244_n8);
   add_244_U7 : OAI21M20D1 port map( A1 => add_244_n7, A2 => a2_in_l_2_port, B 
                           => add_244_n8, Z => add_244_n5);
   add_244_U6 : OAI21D1 port map( A1 => a2_in_l_3_port, A2 => add_244_n5, B => 
                           a2_in_r_3_port, Z => add_244_n6);
   add_244_U5 : OAI21M20D1 port map( A1 => add_244_n5, A2 => a2_in_l_3_port, B 
                           => add_244_n6, Z => add_244_n3);
   add_244_U4 : OAI21D1 port map( A1 => a2_in_l_4_port, A2 => add_244_n3, B => 
                           a2_in_r_4_port, Z => add_244_n4);
   add_244_U3 : OAI21M20D1 port map( A1 => add_244_n3, A2 => a2_in_l_4_port, B 
                           => add_244_n4, Z => add_244_n1);
   add_244_U2 : OAI21D1 port map( A1 => a2_in_l_5_port, A2 => add_244_n1, B => 
                           a2_in_r_5_port, Z => add_244_n2);
   add_244_U1 : OAI21M20D1 port map( A1 => add_244_n1, A2 => a2_in_l_5_port, B 
                           => add_244_n2, Z => add_244_carry_6_port);
   add_244_U1_14 : EXOR3D1 port map( A1 => a2_in_l_14_port, A2 => 
                           a2_in_r_14_port, A3 => add_244_carry_14_port, Z => 
                           N123);
   add_244_U1_6 : ADFULD1 port map( A => a2_in_l_6_port, B => a2_in_r_6_port, 
                           CI => add_244_carry_6_port, CO => 
                           add_244_carry_7_port, S => N115);
   add_244_U1_7 : ADFULD1 port map( A => a2_in_l_7_port, B => a2_in_r_7_port, 
                           CI => add_244_carry_7_port, CO => 
                           add_244_carry_8_port, S => N116);
   add_244_U1_8 : ADFULD1 port map( A => a2_in_l_8_port, B => a2_in_r_8_port, 
                           CI => add_244_carry_8_port, CO => 
                           add_244_carry_9_port, S => N117);
   add_244_U1_9 : ADFULD1 port map( A => a2_in_l_9_port, B => a2_in_r_9_port, 
                           CI => add_244_carry_9_port, CO => 
                           add_244_carry_10_port, S => N118);
   add_244_U1_10 : ADFULD1 port map( A => a2_in_l_10_port, B => a2_in_r_10_port
                           , CI => add_244_carry_10_port, CO => 
                           add_244_carry_11_port, S => N119);
   add_244_U1_11 : ADFULD1 port map( A => a2_in_l_11_port, B => a2_in_r_11_port
                           , CI => add_244_carry_11_port, CO => 
                           add_244_carry_12_port, S => N120);
   add_244_U1_12 : ADFULD1 port map( A => a2_in_l_12_port, B => a2_in_r_12_port
                           , CI => add_244_carry_12_port, CO => 
                           add_244_carry_13_port, S => N121);
   add_244_U1_13 : ADFULD1 port map( A => a2_in_l_13_port, B => a2_in_r_13_port
                           , CI => add_244_carry_13_port, CO => 
                           add_244_carry_14_port, S => N122);
   add_243_U10 : OAI211D1 port map( A1 => a1_in_l_1_port, A2 => a1_in_r_1_port,
                           B => a1_in_l_0_port, C => a1_in_r_0_port, Z => 
                           add_243_n9);
   add_243_U9 : OAI21M20D1 port map( A1 => a1_in_l_1_port, A2 => a1_in_r_1_port
                           , B => add_243_n9, Z => add_243_n7);
   add_243_U8 : OAI21D1 port map( A1 => a1_in_l_2_port, A2 => add_243_n7, B => 
                           a1_in_r_2_port, Z => add_243_n8);
   add_243_U7 : OAI21M20D1 port map( A1 => add_243_n7, A2 => a1_in_l_2_port, B 
                           => add_243_n8, Z => add_243_n5);
   add_243_U6 : OAI21D1 port map( A1 => a1_in_l_3_port, A2 => add_243_n5, B => 
                           a1_in_r_3_port, Z => add_243_n6);
   add_243_U5 : OAI21M20D1 port map( A1 => add_243_n5, A2 => a1_in_l_3_port, B 
                           => add_243_n6, Z => add_243_n3);
   add_243_U4 : OAI21D1 port map( A1 => a1_in_l_4_port, A2 => add_243_n3, B => 
                           a1_in_r_4_port, Z => add_243_n4);
   add_243_U3 : OAI21M20D1 port map( A1 => add_243_n3, A2 => a1_in_l_4_port, B 
                           => add_243_n4, Z => add_243_n1);
   add_243_U2 : OAI21D1 port map( A1 => a1_in_l_5_port, A2 => add_243_n1, B => 
                           a1_in_r_5_port, Z => add_243_n2);
   add_243_U1 : OAI21M20D1 port map( A1 => add_243_n1, A2 => a1_in_l_5_port, B 
                           => add_243_n2, Z => add_243_carry_6_port);
   add_243_U1_14 : EXOR3D1 port map( A1 => a1_in_l_14_port, A2 => 
                           a1_in_r_14_port, A3 => add_243_carry_14_port, Z => 
                           N114);
   add_243_U1_6 : ADFULD1 port map( A => a1_in_l_6_port, B => a1_in_r_6_port, 
                           CI => add_243_carry_6_port, CO => 
                           add_243_carry_7_port, S => N106);
   add_243_U1_7 : ADFULD1 port map( A => a1_in_l_7_port, B => a1_in_r_7_port, 
                           CI => add_243_carry_7_port, CO => 
                           add_243_carry_8_port, S => N107);
   add_243_U1_8 : ADFULD1 port map( A => a1_in_l_8_port, B => a1_in_r_8_port, 
                           CI => add_243_carry_8_port, CO => 
                           add_243_carry_9_port, S => N108);
   add_243_U1_9 : ADFULD1 port map( A => a1_in_l_9_port, B => a1_in_r_9_port, 
                           CI => add_243_carry_9_port, CO => 
                           add_243_carry_10_port, S => N109);
   add_243_U1_10 : ADFULD1 port map( A => a1_in_l_10_port, B => a1_in_r_10_port
                           , CI => add_243_carry_10_port, CO => 
                           add_243_carry_11_port, S => N110);
   add_243_U1_11 : ADFULD1 port map( A => a1_in_l_11_port, B => a1_in_r_11_port
                           , CI => add_243_carry_11_port, CO => 
                           add_243_carry_12_port, S => N111);
   add_243_U1_12 : ADFULD1 port map( A => a1_in_l_12_port, B => a1_in_r_12_port
                           , CI => add_243_carry_12_port, CO => 
                           add_243_carry_13_port, S => N112);
   add_243_U1_13 : ADFULD1 port map( A => a1_in_l_13_port, B => a1_in_r_13_port
                           , CI => add_243_carry_13_port, CO => 
                           add_243_carry_14_port, S => N113);
   mult_238_U121 : NAN2D1 port map( A1 => n193, A2 => m1_in_r_4_port, Z => 
                           mult_238_n23);
   mult_238_U120 : NAN2D1 port map( A1 => n193, A2 => m1_in_r_3_port, Z => 
                           mult_238_n29);
   mult_238_U119 : NAN2D1 port map( A1 => n193, A2 => m1_in_r_2_port, Z => 
                           mult_238_n35);
   mult_238_U118 : NAN2D1 port map( A1 => n193, A2 => m1_in_r_7_port, Z => 
                           mult_238_n46);
   mult_238_U117 : NOR2D1 port map( A1 => mult_238_n121, A2 => mult_238_n119, Z
                           => mult_238_n47);
   mult_238_U116 : NOR2D1 port map( A1 => mult_238_n122, A2 => mult_238_n119, Z
                           => mult_238_n48);
   mult_238_U115 : NOR2D1 port map( A1 => mult_238_n129, A2 => mult_238_n119, Z
                           => mult_238_n49);
   mult_238_U114 : NOR2D1 port map( A1 => mult_238_n130, A2 => mult_238_n119, Z
                           => mult_238_n50);
   mult_238_U113 : NAN2D1 port map( A1 => n193, A2 => m1_in_r_7_port, Z => 
                           mult_238_n51);
   mult_238_U112 : NOR2D1 port map( A1 => mult_238_n121, A2 => mult_238_n119, Z
                           => mult_238_n52);
   mult_238_U111 : NOR2D1 port map( A1 => mult_238_n122, A2 => mult_238_n119, Z
                           => mult_238_n53);
   mult_238_U110 : NOR2D1 port map( A1 => mult_238_n123, A2 => mult_238_n119, Z
                           => mult_238_n54);
   mult_238_U109 : NOR2D1 port map( A1 => mult_238_n125, A2 => mult_238_n119, Z
                           => mult_238_n55);
   mult_238_U108 : NOR2D1 port map( A1 => mult_238_n127, A2 => mult_238_n119, Z
                           => mult_238_n56);
   mult_238_U107 : NOR2D1 port map( A1 => mult_238_n129, A2 => mult_238_n119, Z
                           => mult_238_n57);
   mult_238_U106 : NOR2D1 port map( A1 => mult_238_n130, A2 => mult_238_n119, Z
                           => mult_238_n58);
   mult_238_U105 : NAN2D1 port map( A1 => n193, A2 => m1_in_r_7_port, Z => 
                           mult_238_n59);
   mult_238_U104 : NOR2D1 port map( A1 => mult_238_n121, A2 => mult_238_n119, Z
                           => mult_238_n60);
   mult_238_U103 : NOR2D1 port map( A1 => mult_238_n122, A2 => mult_238_n119, Z
                           => mult_238_n61);
   mult_238_U102 : NOR2D1 port map( A1 => mult_238_n123, A2 => mult_238_n119, Z
                           => mult_238_n62);
   mult_238_U101 : NOR2D1 port map( A1 => mult_238_n125, A2 => mult_238_n119, Z
                           => mult_238_n63);
   mult_238_U100 : NOR2D1 port map( A1 => mult_238_n127, A2 => mult_238_n119, Z
                           => mult_238_n64);
   mult_238_U99 : NOR2D1 port map( A1 => mult_238_n129, A2 => mult_238_n119, Z 
                           => mult_238_n65);
   mult_238_U98 : NOR2D1 port map( A1 => mult_238_n130, A2 => mult_238_n119, Z 
                           => mult_238_n66);
   mult_238_U97 : NAN2D1 port map( A1 => m1_in_r_7_port, A2 => n193, Z => 
                           mult_238_n67);
   mult_238_U96 : NOR2D1 port map( A1 => mult_238_n119, A2 => mult_238_n121, Z 
                           => mult_238_n68);
   mult_238_U95 : NOR2D1 port map( A1 => mult_238_n119, A2 => mult_238_n122, Z 
                           => mult_238_n69);
   mult_238_U94 : NOR2D1 port map( A1 => mult_238_n119, A2 => mult_238_n123, Z 
                           => mult_238_n70);
   mult_238_U93 : NOR2D1 port map( A1 => mult_238_n119, A2 => mult_238_n125, Z 
                           => mult_238_n71);
   mult_238_U92 : NOR2D1 port map( A1 => mult_238_n119, A2 => mult_238_n130, Z 
                           => m1_out_0_port);
   mult_238_U91 : NOR2D1 port map( A1 => mult_238_n119, A2 => mult_238_n129, Z 
                           => m1_out_1_port);
   mult_238_U90 : NOR2D1 port map( A1 => mult_238_n119, A2 => mult_238_n127, Z 
                           => m1_out_2_port);
   mult_238_U89 : INVD1 port map( A => m1_in_r_6_port, Z => mult_238_n121);
   mult_238_U88 : INVD1 port map( A => m1_in_r_5_port, Z => mult_238_n122);
   mult_238_U87 : INVD1 port map( A => m1_in_r_1_port, Z => mult_238_n129);
   mult_238_U86 : INVD1 port map( A => m1_in_r_0_port, Z => mult_238_n130);
   mult_238_U85 : INVD1 port map( A => mult_238_n23, Z => mult_238_n124);
   mult_238_U84 : INVD1 port map( A => mult_238_n29, Z => mult_238_n126);
   mult_238_U83 : INVD1 port map( A => mult_238_n35, Z => mult_238_n128);
   mult_238_U82 : INVD1 port map( A => m1_in_r_2_port, Z => mult_238_n127);
   mult_238_U81 : INVD1 port map( A => m1_in_r_3_port, Z => mult_238_n125);
   mult_238_U80 : INVD1 port map( A => m1_in_r_4_port, Z => mult_238_n123);
   mult_238_U79 : INVD1 port map( A => mult_238_n2, Z => m1_out_15);
   mult_238_U78 : INVD1 port map( A => n193, Z => mult_238_n119);
   mult_238_U30 : ADHALFDL port map( A => mult_238_n65, B => mult_238_n70, CO 
                           => mult_238_n44, S => mult_238_n45);
   mult_238_U29 : ADHALFDL port map( A => mult_238_n50, B => mult_238_n57, CO 
                           => mult_238_n42, S => mult_238_n43);
   mult_238_U28 : ADFULD1 port map( A => mult_238_n64, B => mult_238_n69, CI =>
                           mult_238_n44, CO => mult_238_n40, S => mult_238_n41)
                           ;
   mult_238_U27 : ADFULD1 port map( A => mult_238_n49, B => mult_238_n56, CI =>
                           mult_238_n63, CO => mult_238_n38, S => mult_238_n39)
                           ;
   mult_238_U26 : ADFULD1 port map( A => mult_238_n42, B => mult_238_n68, CI =>
                           mult_238_n39, CO => mult_238_n36, S => mult_238_n37)
                           ;
   mult_238_U24 : ADFULD1 port map( A => mult_238_n55, B => mult_238_n62, CI =>
                           mult_238_n67, CO => mult_238_n32, S => mult_238_n33)
                           ;
   mult_238_U23 : ADFULD1 port map( A => mult_238_n38, B => mult_238_n35, CI =>
                           mult_238_n33, CO => mult_238_n30, S => mult_238_n31)
                           ;
   mult_238_U21 : ADFULD1 port map( A => mult_238_n128, B => mult_238_n61, CI 
                           => mult_238_n54, CO => mult_238_n26, S => 
                           mult_238_n27);
   mult_238_U20 : ADFULD1 port map( A => mult_238_n32, B => mult_238_n29, CI =>
                           mult_238_n27, CO => mult_238_n24, S => mult_238_n25)
                           ;
   mult_238_U18 : ADFULD1 port map( A => mult_238_n126, B => mult_238_n60, CI 
                           => mult_238_n53, CO => mult_238_n20, S => 
                           mult_238_n21);
   mult_238_U17 : ADFULD1 port map( A => mult_238_n26, B => mult_238_n23, CI =>
                           mult_238_n21, CO => mult_238_n18, S => mult_238_n19)
                           ;
   mult_238_U16 : ADFULD1 port map( A => mult_238_n52, B => mult_238_n124, CI 
                           => mult_238_n59, CO => mult_238_n16, S => 
                           mult_238_n17);
   mult_238_U15 : ADFULD1 port map( A => mult_238_n20, B => mult_238_n48, CI =>
                           mult_238_n17, CO => mult_238_n14, S => mult_238_n15)
                           ;
   mult_238_U14 : ADFULD1 port map( A => mult_238_n51, B => mult_238_n47, CI =>
                           mult_238_n16, CO => mult_238_n12, S => mult_238_n13)
                           ;
   mult_238_U13 : ADHALFDL port map( A => mult_238_n71, B => mult_238_n66, CO 
                           => mult_238_n11, S => m1_out_3_port);
   mult_238_U12 : ADFULD1 port map( A => mult_238_n11, B => mult_238_n58, CI =>
                           mult_238_n45, CO => mult_238_n10, S => m1_out_4_port
                           );
   mult_238_U11 : ADFULD1 port map( A => mult_238_n10, B => mult_238_n43, CI =>
                           mult_238_n41, CO => mult_238_n9, S => m1_out_5_port)
                           ;
   mult_238_U10 : ADFULD1 port map( A => mult_238_n37, B => mult_238_n40, CI =>
                           mult_238_n9, CO => mult_238_n8, S => m1_out_6_port);
   mult_238_U9 : ADFULD1 port map( A => mult_238_n31, B => mult_238_n36, CI => 
                           mult_238_n8, CO => mult_238_n7, S => m1_out_7_port);
   mult_238_U8 : ADFULD1 port map( A => mult_238_n25, B => mult_238_n30, CI => 
                           mult_238_n7, CO => mult_238_n6, S => m1_out_8_port);
   mult_238_U7 : ADFULD1 port map( A => mult_238_n19, B => mult_238_n24, CI => 
                           mult_238_n6, CO => mult_238_n5, S => m1_out_9_port);
   mult_238_U6 : ADFULD1 port map( A => mult_238_n15, B => mult_238_n18, CI => 
                           mult_238_n5, CO => mult_238_n4, S => m1_out_10_port)
                           ;
   mult_238_U5 : ADFULD1 port map( A => mult_238_n13, B => mult_238_n14, CI => 
                           mult_238_n4, CO => mult_238_n3, S => m1_out_11_port)
                           ;
   mult_238_U4 : ADFULD1 port map( A => mult_238_n12, B => mult_238_n46, CI => 
                           mult_238_n3, CO => mult_238_n2, S => m1_out_12_port)
                           ;
   mult_242_U121 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m5_in_r_4_port, Z =>
                           mult_242_n23);
   mult_242_U120 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m5_in_r_3_port, Z =>
                           mult_242_n29);
   mult_242_U119 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m5_in_r_2_port, Z =>
                           mult_242_n35);
   mult_242_U118 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m5_in_r_7_port, Z =>
                           mult_242_n46);
   mult_242_U117 : NOR2D1 port map( A1 => mult_242_n121, A2 => mult_242_n119, Z
                           => mult_242_n47);
   mult_242_U116 : NOR2D1 port map( A1 => mult_242_n122, A2 => mult_242_n119, Z
                           => mult_242_n48);
   mult_242_U115 : NOR2D1 port map( A1 => mult_242_n129, A2 => mult_242_n119, Z
                           => mult_242_n49);
   mult_242_U114 : NOR2D1 port map( A1 => mult_242_n130, A2 => mult_242_n119, Z
                           => mult_242_n50);
   mult_242_U113 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m5_in_r_7_port, Z =>
                           mult_242_n51);
   mult_242_U112 : NOR2D1 port map( A1 => mult_242_n121, A2 => mult_242_n119, Z
                           => mult_242_n52);
   mult_242_U111 : NOR2D1 port map( A1 => mult_242_n122, A2 => mult_242_n119, Z
                           => mult_242_n53);
   mult_242_U110 : NOR2D1 port map( A1 => mult_242_n123, A2 => mult_242_n119, Z
                           => mult_242_n54);
   mult_242_U109 : NOR2D1 port map( A1 => mult_242_n125, A2 => mult_242_n119, Z
                           => mult_242_n55);
   mult_242_U108 : NOR2D1 port map( A1 => mult_242_n127, A2 => mult_242_n119, Z
                           => mult_242_n56);
   mult_242_U107 : NOR2D1 port map( A1 => mult_242_n129, A2 => mult_242_n119, Z
                           => mult_242_n57);
   mult_242_U106 : NOR2D1 port map( A1 => mult_242_n130, A2 => mult_242_n119, Z
                           => mult_242_n58);
   mult_242_U105 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m5_in_r_7_port, Z =>
                           mult_242_n59);
   mult_242_U104 : NOR2D1 port map( A1 => mult_242_n121, A2 => mult_242_n119, Z
                           => mult_242_n60);
   mult_242_U103 : NOR2D1 port map( A1 => mult_242_n122, A2 => mult_242_n119, Z
                           => mult_242_n61);
   mult_242_U102 : NOR2D1 port map( A1 => mult_242_n123, A2 => mult_242_n119, Z
                           => mult_242_n62);
   mult_242_U101 : NOR2D1 port map( A1 => mult_242_n125, A2 => mult_242_n119, Z
                           => mult_242_n63);
   mult_242_U100 : NOR2D1 port map( A1 => mult_242_n127, A2 => mult_242_n119, Z
                           => mult_242_n64);
   mult_242_U99 : NOR2D1 port map( A1 => mult_242_n129, A2 => mult_242_n119, Z 
                           => mult_242_n65);
   mult_242_U98 : NOR2D1 port map( A1 => mult_242_n130, A2 => mult_242_n119, Z 
                           => mult_242_n66);
   mult_242_U97 : NAN2D1 port map( A1 => m5_in_r_7_port, A2 => m5_in_l_0, Z => 
                           mult_242_n67);
   mult_242_U96 : NOR2D1 port map( A1 => mult_242_n119, A2 => mult_242_n121, Z 
                           => mult_242_n68);
   mult_242_U95 : NOR2D1 port map( A1 => mult_242_n119, A2 => mult_242_n122, Z 
                           => mult_242_n69);
   mult_242_U94 : NOR2D1 port map( A1 => mult_242_n119, A2 => mult_242_n123, Z 
                           => mult_242_n70);
   mult_242_U93 : NOR2D1 port map( A1 => mult_242_n119, A2 => mult_242_n125, Z 
                           => mult_242_n71);
   mult_242_U92 : NOR2D1 port map( A1 => mult_242_n119, A2 => mult_242_n130, Z 
                           => m5_out_0_port);
   mult_242_U91 : NOR2D1 port map( A1 => mult_242_n119, A2 => mult_242_n129, Z 
                           => m5_out_1_port);
   mult_242_U90 : NOR2D1 port map( A1 => mult_242_n119, A2 => mult_242_n127, Z 
                           => m5_out_2_port);
   mult_242_U89 : INVD1 port map( A => m5_in_r_6_port, Z => mult_242_n121);
   mult_242_U88 : INVD1 port map( A => m5_in_r_5_port, Z => mult_242_n122);
   mult_242_U87 : INVD1 port map( A => m5_in_r_0_port, Z => mult_242_n130);
   mult_242_U86 : INVD1 port map( A => m5_in_r_1_port, Z => mult_242_n129);
   mult_242_U85 : INVD1 port map( A => mult_242_n23, Z => mult_242_n124);
   mult_242_U84 : INVD1 port map( A => mult_242_n29, Z => mult_242_n126);
   mult_242_U83 : INVD1 port map( A => mult_242_n35, Z => mult_242_n128);
   mult_242_U82 : INVD1 port map( A => m5_in_r_3_port, Z => mult_242_n125);
   mult_242_U81 : INVD1 port map( A => m5_in_r_2_port, Z => mult_242_n127);
   mult_242_U80 : INVD1 port map( A => m5_in_r_4_port, Z => mult_242_n123);
   mult_242_U79 : INVD1 port map( A => mult_242_n2, Z => m5_out_15);
   mult_242_U78 : INVD1 port map( A => m5_in_l_0, Z => mult_242_n119);
   mult_242_U30 : ADHALFDL port map( A => mult_242_n65, B => mult_242_n70, CO 
                           => mult_242_n44, S => mult_242_n45);
   mult_242_U29 : ADHALFDL port map( A => mult_242_n50, B => mult_242_n57, CO 
                           => mult_242_n42, S => mult_242_n43);
   mult_242_U28 : ADFULD1 port map( A => mult_242_n64, B => mult_242_n69, CI =>
                           mult_242_n44, CO => mult_242_n40, S => mult_242_n41)
                           ;
   mult_242_U27 : ADFULD1 port map( A => mult_242_n49, B => mult_242_n56, CI =>
                           mult_242_n63, CO => mult_242_n38, S => mult_242_n39)
                           ;
   mult_242_U26 : ADFULD1 port map( A => mult_242_n42, B => mult_242_n68, CI =>
                           mult_242_n39, CO => mult_242_n36, S => mult_242_n37)
                           ;
   mult_242_U24 : ADFULD1 port map( A => mult_242_n55, B => mult_242_n62, CI =>
                           mult_242_n67, CO => mult_242_n32, S => mult_242_n33)
                           ;
   mult_242_U23 : ADFULD1 port map( A => mult_242_n38, B => mult_242_n35, CI =>
                           mult_242_n33, CO => mult_242_n30, S => mult_242_n31)
                           ;
   mult_242_U21 : ADFULD1 port map( A => mult_242_n128, B => mult_242_n61, CI 
                           => mult_242_n54, CO => mult_242_n26, S => 
                           mult_242_n27);
   mult_242_U20 : ADFULD1 port map( A => mult_242_n32, B => mult_242_n29, CI =>
                           mult_242_n27, CO => mult_242_n24, S => mult_242_n25)
                           ;
   mult_242_U18 : ADFULD1 port map( A => mult_242_n126, B => mult_242_n60, CI 
                           => mult_242_n53, CO => mult_242_n20, S => 
                           mult_242_n21);
   mult_242_U17 : ADFULD1 port map( A => mult_242_n26, B => mult_242_n23, CI =>
                           mult_242_n21, CO => mult_242_n18, S => mult_242_n19)
                           ;
   mult_242_U16 : ADFULD1 port map( A => mult_242_n52, B => mult_242_n124, CI 
                           => mult_242_n59, CO => mult_242_n16, S => 
                           mult_242_n17);
   mult_242_U15 : ADFULD1 port map( A => mult_242_n20, B => mult_242_n48, CI =>
                           mult_242_n17, CO => mult_242_n14, S => mult_242_n15)
                           ;
   mult_242_U14 : ADFULD1 port map( A => mult_242_n51, B => mult_242_n47, CI =>
                           mult_242_n16, CO => mult_242_n12, S => mult_242_n13)
                           ;
   mult_242_U13 : ADHALFDL port map( A => mult_242_n71, B => mult_242_n66, CO 
                           => mult_242_n11, S => m5_out_3_port);
   mult_242_U12 : ADFULD1 port map( A => mult_242_n11, B => mult_242_n58, CI =>
                           mult_242_n45, CO => mult_242_n10, S => m5_out_4_port
                           );
   mult_242_U11 : ADFULD1 port map( A => mult_242_n10, B => mult_242_n43, CI =>
                           mult_242_n41, CO => mult_242_n9, S => m5_out_5_port)
                           ;
   mult_242_U10 : ADFULD1 port map( A => mult_242_n37, B => mult_242_n40, CI =>
                           mult_242_n9, CO => mult_242_n8, S => m5_out_6_port);
   mult_242_U9 : ADFULD1 port map( A => mult_242_n31, B => mult_242_n36, CI => 
                           mult_242_n8, CO => mult_242_n7, S => m5_out_7_port);
   mult_242_U8 : ADFULD1 port map( A => mult_242_n25, B => mult_242_n30, CI => 
                           mult_242_n7, CO => mult_242_n6, S => m5_out_8_port);
   mult_242_U7 : ADFULD1 port map( A => mult_242_n19, B => mult_242_n24, CI => 
                           mult_242_n6, CO => mult_242_n5, S => m5_out_9_port);
   mult_242_U6 : ADFULD1 port map( A => mult_242_n15, B => mult_242_n18, CI => 
                           mult_242_n5, CO => mult_242_n4, S => m5_out_10_port)
                           ;
   mult_242_U5 : ADFULD1 port map( A => mult_242_n13, B => mult_242_n14, CI => 
                           mult_242_n4, CO => mult_242_n3, S => m5_out_11_port)
                           ;
   mult_242_U4 : ADFULD1 port map( A => mult_242_n12, B => mult_242_n46, CI => 
                           mult_242_n3, CO => mult_242_n2, S => m5_out_12_port)
                           ;
   mult_240_U121 : AND2D1 port map( A1 => m4_in_r_6_port, A2 => m5_in_l_0, Z =>
                           mult_240_n14);
   mult_240_U120 : NAN2D1 port map( A1 => m4_in_r_5_port, A2 => m5_in_l_0, Z =>
                           mult_240_n15);
   mult_240_U119 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_6_port, Z =>
                           mult_240_n28);
   mult_240_U118 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_4_port, Z =>
                           mult_240_n34);
   mult_240_U117 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_4_port, Z =>
                           mult_240_n129);
   mult_240_U116 : NAN2D1 port map( A1 => m4_in_r_6_port, A2 => m5_in_l_0, Z =>
                           mult_240_n130);
   mult_240_U115 : NAN2D1 port map( A1 => mult_240_n129, A2 => mult_240_n130, Z
                           => mult_240_n37);
   mult_240_U114 : EXNOR2D1 port map( A1 => mult_240_n129, A2 => mult_240_n130,
                           Z => mult_240_n38);
   mult_240_U113 : NAN2D1 port map( A1 => m4_in_r_4_port, A2 => m5_in_l_0, Z =>
                           mult_240_n46);
   mult_240_U112 : NAN2D1 port map( A1 => m4_in_r_3_port, A2 => m5_in_l_0, Z =>
                           mult_240_n47);
   mult_240_U111 : NAN2D1 port map( A1 => m4_in_r_2_port, A2 => m5_in_l_0, Z =>
                           mult_240_n48);
   mult_240_U110 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_1_port, Z =>
                           mult_240_n49);
   mult_240_U109 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_0_port, Z =>
                           mult_240_n50);
   mult_240_U108 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z =>
                           mult_240_n51);
   mult_240_U107 : NOR2M1D1 port map( A1 => m4_in_r_6_port, A2 => mult_240_n119
                           , Z => mult_240_n52);
   mult_240_U106 : NOR2D1 port map( A1 => mult_240_n121, A2 => mult_240_n119, Z
                           => mult_240_n53);
   mult_240_U105 : NOR2D1 port map( A1 => mult_240_n124, A2 => mult_240_n119, Z
                           => mult_240_n54);
   mult_240_U104 : NOR2D1 port map( A1 => mult_240_n125, A2 => mult_240_n119, Z
                           => mult_240_n55);
   mult_240_U103 : NOR2D1 port map( A1 => mult_240_n126, A2 => mult_240_n119, Z
                           => mult_240_n56);
   mult_240_U102 : NOR2D1 port map( A1 => mult_240_n127, A2 => mult_240_n119, Z
                           => mult_240_n57);
   mult_240_U101 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z =>
                           mult_240_n58);
   mult_240_U100 : NOR2D1 port map( A1 => mult_240_n121, A2 => mult_240_n119, Z
                           => mult_240_n59);
   mult_240_U99 : NOR2D1 port map( A1 => mult_240_n124, A2 => mult_240_n119, Z 
                           => mult_240_n61);
   mult_240_U98 : NOR2D1 port map( A1 => mult_240_n125, A2 => mult_240_n119, Z 
                           => mult_240_n62);
   mult_240_U97 : NOR2D1 port map( A1 => mult_240_n126, A2 => mult_240_n119, Z 
                           => mult_240_n63);
   mult_240_U96 : NOR2D1 port map( A1 => mult_240_n127, A2 => mult_240_n119, Z 
                           => mult_240_n64);
   mult_240_U95 : NAN2D1 port map( A1 => m4_in_r_7_port, A2 => m5_in_l_0, Z => 
                           mult_240_n65);
   mult_240_U94 : NOR2D1 port map( A1 => mult_240_n119, A2 => mult_240_n121, Z 
                           => mult_240_n67);
   mult_240_U93 : NOR2M1D1 port map( A1 => m4_in_r_4_port, A2 => mult_240_n119,
                           Z => mult_240_n68);
   mult_240_U92 : NOR2D1 port map( A1 => mult_240_n119, A2 => mult_240_n124, Z 
                           => mult_240_n69);
   mult_240_U91 : NOR2D1 port map( A1 => mult_240_n119, A2 => mult_240_n125, Z 
                           => mult_240_n70);
   mult_240_U90 : AND2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z => 
                           mult_240_n128);
   mult_240_U89 : EXNOR3D1 port map( A1 => mult_240_n2, A2 => mult_240_n128, A3
                           => mult_240_n14, Z => m3_out_14_port);
   mult_240_U88 : NOR2D1 port map( A1 => mult_240_n119, A2 => mult_240_n127, Z 
                           => m3_out_1_port);
   mult_240_U87 : NOR2D1 port map( A1 => mult_240_n119, A2 => mult_240_n126, Z 
                           => m3_out_2_port);
   mult_240_U86 : INVD1 port map( A => mult_240_n28, Z => mult_240_n120);
   mult_240_U85 : INVD1 port map( A => mult_240_n34, Z => mult_240_n123);
   mult_240_U84 : INVD1 port map( A => m4_in_r_5_port, Z => mult_240_n121);
   mult_240_U83 : INVD1 port map( A => m4_in_r_0_port, Z => mult_240_n127);
   mult_240_U82 : INVD1 port map( A => m4_in_r_2_port, Z => mult_240_n125);
   mult_240_U81 : INVD1 port map( A => m4_in_r_1_port, Z => mult_240_n126);
   mult_240_U80 : INVD1 port map( A => m4_in_r_3_port, Z => mult_240_n124);
   mult_240_U79 : INVD1 port map( A => mult_240_n15, Z => mult_240_n122);
   mult_240_U78 : INVD1 port map( A => m5_in_l_0, Z => mult_240_n119);
   mult_240_U30 : ADHALFDL port map( A => mult_240_n63, B => mult_240_n69, CO 
                           => mult_240_n43, S => mult_240_n44);
   mult_240_U29 : ADFULD1 port map( A => mult_240_n56, B => mult_240_n68, CI =>
                           mult_240_n62, CO => mult_240_n41, S => mult_240_n42)
                           ;
   mult_240_U28 : ADFULD1 port map( A => mult_240_n55, B => mult_240_n67, CI =>
                           mult_240_n61, CO => mult_240_n39, S => mult_240_n40)
                           ;
   mult_240_U25 : ADFULD1 port map( A => mult_240_n50, B => mult_240_n54, CI =>
                           mult_240_n38, CO => mult_240_n35, S => mult_240_n36)
                           ;
   mult_240_U23 : ADFULD1 port map( A => mult_240_n65, B => mult_240_n59, CI =>
                           mult_240_n49, CO => mult_240_n31, S => mult_240_n32)
                           ;
   mult_240_U22 : ADFULD1 port map( A => mult_240_n37, B => mult_240_n34, CI =>
                           mult_240_n32, CO => mult_240_n29, S => mult_240_n30)
                           ;
   mult_240_U20 : ADFULD1 port map( A => mult_240_n123, B => mult_240_n53, CI 
                           => mult_240_n48, CO => mult_240_n25, S => 
                           mult_240_n26);
   mult_240_U19 : ADFULD1 port map( A => mult_240_n31, B => mult_240_n28, CI =>
                           mult_240_n26, CO => mult_240_n23, S => mult_240_n24)
                           ;
   mult_240_U18 : ADFULD1 port map( A => mult_240_n52, B => mult_240_n120, CI 
                           => mult_240_n47, CO => mult_240_n21, S => 
                           mult_240_n22);
   mult_240_U17 : ADFULD1 port map( A => mult_240_n25, B => mult_240_n58, CI =>
                           mult_240_n22, CO => mult_240_n19, S => mult_240_n20)
                           ;
   mult_240_U16 : ADFULD1 port map( A => mult_240_n46, B => mult_240_n51, CI =>
                           mult_240_n21, CO => mult_240_n17, S => mult_240_n18)
                           ;
   mult_240_U13 : ADHALFDL port map( A => mult_240_n70, B => mult_240_n64, CO 
                           => mult_240_n12, S => m3_out_3_port);
   mult_240_U12 : ADFULD1 port map( A => mult_240_n12, B => mult_240_n57, CI =>
                           mult_240_n44, CO => mult_240_n11, S => m3_out_4_port
                           );
   mult_240_U11 : ADFULD1 port map( A => mult_240_n42, B => mult_240_n43, CI =>
                           mult_240_n11, CO => mult_240_n10, S => m3_out_5_port
                           );
   mult_240_U10 : ADFULD1 port map( A => mult_240_n40, B => mult_240_n41, CI =>
                           mult_240_n10, CO => mult_240_n9, S => m3_out_6_port)
                           ;
   mult_240_U9 : ADFULD1 port map( A => mult_240_n36, B => mult_240_n39, CI => 
                           mult_240_n9, CO => mult_240_n8, S => m3_out_7_port);
   mult_240_U8 : ADFULD1 port map( A => mult_240_n30, B => mult_240_n35, CI => 
                           mult_240_n8, CO => mult_240_n7, S => m3_out_8_port);
   mult_240_U7 : ADFULD1 port map( A => mult_240_n24, B => mult_240_n29, CI => 
                           mult_240_n7, CO => mult_240_n6, S => m3_out_9_port);
   mult_240_U6 : ADFULD1 port map( A => mult_240_n20, B => mult_240_n23, CI => 
                           mult_240_n6, CO => mult_240_n5, S => m3_out_10_port)
                           ;
   mult_240_U5 : ADFULD1 port map( A => mult_240_n18, B => mult_240_n19, CI => 
                           mult_240_n5, CO => mult_240_n4, S => m3_out_11_port)
                           ;
   mult_240_U4 : ADFULD1 port map( A => mult_240_n17, B => mult_240_n122, CI =>
                           mult_240_n4, CO => mult_240_n3, S => m3_out_12_port)
                           ;
   mult_240_U3 : ADFULD1 port map( A => mult_240_n14, B => mult_240_n15, CI => 
                           mult_240_n3, CO => mult_240_n2, S => m3_out_13_port)
                           ;
   mult_241_U170 : NOR2D1 port map( A1 => mult_241_n176, A2 => mult_241_n167, Z
                           => mult_241_n100);
   mult_241_U169 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z =>
                           mult_241_n101);
   mult_241_U168 : NOR2D1 port map( A1 => mult_241_n169, A2 => mult_241_n167, Z
                           => mult_241_n102);
   mult_241_U167 : NOR2D1 port map( A1 => mult_241_n171, A2 => mult_241_n167, Z
                           => mult_241_n103);
   mult_241_U166 : NOR2D1 port map( A1 => mult_241_n172, A2 => mult_241_n167, Z
                           => mult_241_n104);
   mult_241_U165 : NOR2D1 port map( A1 => mult_241_n173, A2 => mult_241_n167, Z
                           => mult_241_n105);
   mult_241_U164 : NOR2D1 port map( A1 => mult_241_n174, A2 => mult_241_n167, Z
                           => mult_241_n106);
   mult_241_U163 : NOR2D1 port map( A1 => mult_241_n175, A2 => mult_241_n167, Z
                           => mult_241_n107);
   mult_241_U162 : NOR2D1 port map( A1 => mult_241_n176, A2 => mult_241_n167, Z
                           => mult_241_n108);
   mult_241_U161 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z =>
                           mult_241_n109);
   mult_241_U160 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n169, Z
                           => mult_241_n110);
   mult_241_U159 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n171, Z
                           => mult_241_n111);
   mult_241_U158 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n172, Z
                           => mult_241_n112);
   mult_241_U157 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n173, Z
                           => mult_241_n113);
   mult_241_U156 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n174, Z
                           => mult_241_n114);
   mult_241_U155 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n175, Z
                           => mult_241_n115);
   mult_241_U154 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_6_port, Z =>
                           mult_241_n20);
   mult_241_U153 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_5_port, Z =>
                           mult_241_n24);
   mult_241_U152 : NAN2D1 port map( A1 => m4_in_r_6_port, A2 => m5_in_l_0, Z =>
                           mult_241_n179);
   mult_241_U151 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_2_port, Z =>
                           mult_241_n178);
   mult_241_U150 : NAN2D1 port map( A1 => mult_241_n179, A2 => mult_241_n178, Z
                           => mult_241_n41);
   mult_241_U149 : EXNOR2D1 port map( A1 => mult_241_n178, A2 => mult_241_n179,
                           Z => mult_241_n42);
   mult_241_U148 : NAN2D1 port map( A1 => m4_in_r_6_port, A2 => m5_in_l_0, Z =>
                           mult_241_n72);
   mult_241_U147 : NAN2D1 port map( A1 => m4_in_r_5_port, A2 => m5_in_l_0, Z =>
                           mult_241_n73);
   mult_241_U146 : NAN2D1 port map( A1 => m4_in_r_4_port, A2 => m5_in_l_0, Z =>
                           mult_241_n74);
   mult_241_U145 : NAN2D1 port map( A1 => m4_in_r_3_port, A2 => m5_in_l_0, Z =>
                           mult_241_n75);
   mult_241_U144 : NAN2D1 port map( A1 => m4_in_r_2_port, A2 => m5_in_l_0, Z =>
                           mult_241_n76);
   mult_241_U143 : NAN2D1 port map( A1 => m4_in_r_1_port, A2 => m5_in_l_0, Z =>
                           mult_241_n77);
   mult_241_U142 : NAN2D1 port map( A1 => m4_in_r_0_port, A2 => m5_in_l_0, Z =>
                           mult_241_n78);
   mult_241_U141 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z =>
                           mult_241_n79);
   mult_241_U140 : NOR2D1 port map( A1 => mult_241_n172, A2 => mult_241_n167, Z
                           => mult_241_n80);
   mult_241_U139 : NOR2D1 port map( A1 => mult_241_n173, A2 => mult_241_n167, Z
                           => mult_241_n81);
   mult_241_U138 : NOR2D1 port map( A1 => mult_241_n175, A2 => mult_241_n167, Z
                           => mult_241_n83);
   mult_241_U137 : NOR2D1 port map( A1 => mult_241_n176, A2 => mult_241_n167, Z
                           => mult_241_n84);
   mult_241_U136 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z =>
                           mult_241_n85);
   mult_241_U135 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n169, Z
                           => mult_241_n86);
   mult_241_U134 : NOR2D1 port map( A1 => mult_241_n171, A2 => mult_241_n167, Z
                           => mult_241_n87);
   mult_241_U133 : NOR2D1 port map( A1 => mult_241_n172, A2 => mult_241_n167, Z
                           => mult_241_n88);
   mult_241_U132 : NOR2D1 port map( A1 => mult_241_n173, A2 => mult_241_n167, Z
                           => mult_241_n89);
   mult_241_U131 : NOR2D1 port map( A1 => mult_241_n174, A2 => mult_241_n167, Z
                           => mult_241_n90);
   mult_241_U130 : NOR2D1 port map( A1 => mult_241_n175, A2 => mult_241_n167, Z
                           => mult_241_n91);
   mult_241_U129 : NOR2D1 port map( A1 => mult_241_n176, A2 => mult_241_n167, Z
                           => mult_241_n92);
   mult_241_U128 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z =>
                           mult_241_n93);
   mult_241_U127 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n171, Z
                           => mult_241_n95);
   mult_241_U126 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n172, Z
                           => mult_241_n96);
   mult_241_U125 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n173, Z
                           => mult_241_n97);
   mult_241_U124 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n174, Z
                           => mult_241_n98);
   mult_241_U123 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n175, Z
                           => mult_241_n99);
   mult_241_U122 : NOR2D1 port map( A1 => mult_241_n167, A2 => mult_241_n176, Z
                           => m4_out_0_port);
   mult_241_U121 : AND2D1 port map( A1 => m5_in_l_0, A2 => m4_in_r_7_port, Z =>
                           mult_241_n177);
   mult_241_U120 : EXOR3D1 port map( A1 => mult_241_n2, A2 => mult_241_n15, A3 
                           => mult_241_n177, Z => m4_out_14_port);
   mult_241_U119 : INVD1 port map( A => mult_241_n20, Z => mult_241_n168);
   mult_241_U118 : INVD1 port map( A => mult_241_n24, Z => mult_241_n170);
   mult_241_U117 : INVD1 port map( A => m4_in_r_5_port, Z => mult_241_n171);
   mult_241_U116 : INVD1 port map( A => m4_in_r_6_port, Z => mult_241_n169);
   mult_241_U115 : INVD1 port map( A => m4_in_r_4_port, Z => mult_241_n172);
   mult_241_U114 : INVD1 port map( A => m4_in_r_0_port, Z => mult_241_n176);
   mult_241_U113 : INVD1 port map( A => m4_in_r_3_port, Z => mult_241_n173);
   mult_241_U112 : INVD1 port map( A => m4_in_r_1_port, Z => mult_241_n175);
   mult_241_U111 : INVD1 port map( A => m4_in_r_2_port, Z => mult_241_n174);
   mult_241_U110 : INVD1 port map( A => m5_in_l_0, Z => mult_241_n167);
   mult_241_U44 : ADHALFDL port map( A => mult_241_n107, B => mult_241_n114, CO
                           => mult_241_n69, S => mult_241_n70);
   mult_241_U43 : ADHALFDL port map( A => mult_241_n92, B => mult_241_n99, CO 
                           => mult_241_n67, S => mult_241_n68);
   mult_241_U42 : ADFULD1 port map( A => mult_241_n106, B => mult_241_n113, CI 
                           => mult_241_n69, CO => mult_241_n65, S => 
                           mult_241_n66);
   mult_241_U41 : ADFULD1 port map( A => mult_241_n91, B => mult_241_n98, CI =>
                           mult_241_n105, CO => mult_241_n63, S => mult_241_n64
                           );
   mult_241_U40 : ADFULD1 port map( A => mult_241_n67, B => mult_241_n112, CI 
                           => mult_241_n64, CO => mult_241_n61, S => 
                           mult_241_n62);
   mult_241_U39 : ADFULD1 port map( A => mult_241_n90, B => mult_241_n97, CI =>
                           mult_241_n104, CO => mult_241_n59, S => mult_241_n60
                           );
   mult_241_U38 : ADFULD1 port map( A => mult_241_n63, B => mult_241_n111, CI 
                           => mult_241_n60, CO => mult_241_n57, S => 
                           mult_241_n58);
   mult_241_U37 : ADHALFDL port map( A => mult_241_n84, B => mult_241_n89, CO 
                           => mult_241_n55, S => mult_241_n56);
   mult_241_U36 : ADFULD1 port map( A => mult_241_n96, B => mult_241_n110, CI 
                           => mult_241_n103, CO => mult_241_n53, S => 
                           mult_241_n54);
   mult_241_U35 : ADFULD1 port map( A => mult_241_n59, B => mult_241_n56, CI =>
                           mult_241_n54, CO => mult_241_n51, S => mult_241_n52)
                           ;
   mult_241_U34 : ADHALFDL port map( A => mult_241_n95, B => mult_241_n88, CO 
                           => mult_241_n49, S => mult_241_n50);
   mult_241_U33 : ADFULD1 port map( A => mult_241_n83, B => mult_241_n102, CI 
                           => mult_241_n78, CO => mult_241_n47, S => 
                           mult_241_n48);
   mult_241_U32 : ADFULD1 port map( A => mult_241_n55, B => mult_241_n109, CI 
                           => mult_241_n50, CO => mult_241_n45, S => 
                           mult_241_n46);
   mult_241_U31 : ADFULD1 port map( A => mult_241_n48, B => mult_241_n53, CI =>
                           mult_241_n46, CO => mult_241_n43, S => mult_241_n44)
                           ;
   mult_241_U28 : ADFULD1 port map( A => mult_241_n101, B => mult_241_n87, CI 
                           => mult_241_n77, CO => mult_241_n39, S => 
                           mult_241_n40);
   mult_241_U27 : ADFULD1 port map( A => mult_241_n42, B => mult_241_n49, CI =>
                           mult_241_n47, CO => mult_241_n37, S => mult_241_n38)
                           ;
   mult_241_U26 : ADFULD1 port map( A => mult_241_n45, B => mult_241_n40, CI =>
                           mult_241_n38, CO => mult_241_n35, S => mult_241_n36)
                           ;
   mult_241_U25 : ADFULD1 port map( A => mult_241_n81, B => mult_241_n86, CI =>
                           mult_241_n76, CO => mult_241_n33, S => mult_241_n34)
                           ;
   mult_241_U24 : ADFULD1 port map( A => mult_241_n41, B => mult_241_n93, CI =>
                           mult_241_n39, CO => mult_241_n31, S => mult_241_n32)
                           ;
   mult_241_U23 : ADFULD1 port map( A => mult_241_n37, B => mult_241_n34, CI =>
                           mult_241_n32, CO => mult_241_n29, S => mult_241_n30)
                           ;
   mult_241_U22 : ADFULD1 port map( A => mult_241_n85, B => mult_241_n80, CI =>
                           mult_241_n75, CO => mult_241_n27, S => mult_241_n28)
                           ;
   mult_241_U21 : ADFULD1 port map( A => mult_241_n28, B => mult_241_n33, CI =>
                           mult_241_n31, CO => mult_241_n25, S => mult_241_n26)
                           ;
   mult_241_U19 : ADFULD1 port map( A => mult_241_n24, B => mult_241_n74, CI =>
                           mult_241_n27, CO => mult_241_n21, S => mult_241_n22)
                           ;
   mult_241_U17 : ADFULD1 port map( A => mult_241_n73, B => mult_241_n170, CI 
                           => mult_241_n20, CO => mult_241_n17, S => 
                           mult_241_n18);
   mult_241_U16 : ADFULD1 port map( A => mult_241_n79, B => mult_241_n168, CI 
                           => mult_241_n72, CO => mult_241_n15, S => 
                           mult_241_n16);
   mult_241_U15 : ADHALFDL port map( A => mult_241_n115, B => mult_241_n108, CO
                           => mult_241_n14, S => m4_out_1_port);
   mult_241_U14 : ADFULD1 port map( A => mult_241_n14, B => mult_241_n100, CI 
                           => mult_241_n70, CO => mult_241_n13, S => 
                           m4_out_2_port);
   mult_241_U13 : ADFULD1 port map( A => mult_241_n13, B => mult_241_n68, CI =>
                           mult_241_n66, CO => mult_241_n12, S => m4_out_3_port
                           );
   mult_241_U12 : ADFULD1 port map( A => mult_241_n62, B => mult_241_n65, CI =>
                           mult_241_n12, CO => mult_241_n11, S => m4_out_4_port
                           );
   mult_241_U11 : ADFULD1 port map( A => mult_241_n58, B => mult_241_n61, CI =>
                           mult_241_n11, CO => mult_241_n10, S => m4_out_5_port
                           );
   mult_241_U10 : ADFULD1 port map( A => mult_241_n52, B => mult_241_n57, CI =>
                           mult_241_n10, CO => mult_241_n9, S => m4_out_6_port)
                           ;
   mult_241_U9 : ADFULD1 port map( A => mult_241_n44, B => mult_241_n51, CI => 
                           mult_241_n9, CO => mult_241_n8, S => m4_out_7_port);
   mult_241_U8 : ADFULD1 port map( A => mult_241_n36, B => mult_241_n43, CI => 
                           mult_241_n8, CO => mult_241_n7, S => m4_out_8_port);
   mult_241_U7 : ADFULD1 port map( A => mult_241_n30, B => mult_241_n35, CI => 
                           mult_241_n7, CO => mult_241_n6, S => m4_out_9_port);
   mult_241_U6 : ADFULD1 port map( A => mult_241_n26, B => mult_241_n29, CI => 
                           mult_241_n6, CO => mult_241_n5, S => m4_out_10_port)
                           ;
   mult_241_U5 : ADFULD1 port map( A => mult_241_n25, B => mult_241_n22, CI => 
                           mult_241_n5, CO => mult_241_n4, S => m4_out_11_port)
                           ;
   mult_241_U4 : ADFULD1 port map( A => mult_241_n21, B => mult_241_n18, CI => 
                           mult_241_n4, CO => mult_241_n3, S => m4_out_12_port)
                           ;
   mult_241_U3 : ADFULD1 port map( A => mult_241_n16, B => mult_241_n17, CI => 
                           mult_241_n3, CO => mult_241_n2, S => m4_out_13_port)
                           ;
   mult_239_U98 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m2_in_r_6_port, Z => 
                           mult_239_n15);
   mult_239_U97 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m2_in_r_5_port, Z => 
                           mult_239_n17);
   mult_239_U96 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m2_in_r_4_port, Z => 
                           mult_239_n19);
   mult_239_U95 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m2_in_r_3_port, Z => 
                           mult_239_n21);
   mult_239_U94 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m2_in_r_1_port, Z => 
                           mult_239_n27);
   mult_239_U93 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m2_in_r_7_port, Z => 
                           mult_239_n30);
   mult_239_U92 : NOR2D1 port map( A1 => mult_239_n106, A2 => mult_239_n96, Z 
                           => mult_239_n31);
   mult_239_U91 : NOR2D1 port map( A1 => mult_239_n109, A2 => mult_239_n96, Z 
                           => mult_239_n32);
   mult_239_U90 : NAN2D1 port map( A1 => m5_in_l_0, A2 => m2_in_r_7_port, Z => 
                           mult_239_n33);
   mult_239_U89 : NOR2D1 port map( A1 => mult_239_n98, A2 => mult_239_n96, Z =>
                           mult_239_n34);
   mult_239_U88 : NOR2D1 port map( A1 => mult_239_n100, A2 => mult_239_n96, Z 
                           => mult_239_n35);
   mult_239_U87 : NOR2D1 port map( A1 => mult_239_n102, A2 => mult_239_n96, Z 
                           => mult_239_n36);
   mult_239_U86 : NOR2D1 port map( A1 => mult_239_n104, A2 => mult_239_n96, Z 
                           => mult_239_n37);
   mult_239_U85 : NOR2D1 port map( A1 => mult_239_n106, A2 => mult_239_n96, Z 
                           => mult_239_n38);
   mult_239_U84 : NOR2D1 port map( A1 => mult_239_n107, A2 => mult_239_n96, Z 
                           => mult_239_n39);
   mult_239_U83 : NOR2D1 port map( A1 => mult_239_n109, A2 => mult_239_n96, Z 
                           => mult_239_n40);
   mult_239_U82 : NAN2D1 port map( A1 => m2_in_r_7_port, A2 => m5_in_l_0, Z => 
                           mult_239_n41);
   mult_239_U81 : NOR2D1 port map( A1 => mult_239_n96, A2 => mult_239_n98, Z =>
                           mult_239_n42);
   mult_239_U80 : NOR2D1 port map( A1 => mult_239_n96, A2 => mult_239_n100, Z 
                           => mult_239_n43);
   mult_239_U79 : NOR2D1 port map( A1 => mult_239_n96, A2 => mult_239_n102, Z 
                           => mult_239_n44);
   mult_239_U78 : NOR2D1 port map( A1 => mult_239_n96, A2 => mult_239_n104, Z 
                           => mult_239_n45);
   mult_239_U77 : NOR2D1 port map( A1 => mult_239_n96, A2 => mult_239_n106, Z 
                           => mult_239_n46);
   mult_239_U76 : NOR2D1 port map( A1 => mult_239_n96, A2 => mult_239_n107, Z 
                           => mult_239_n47);
   mult_239_U75 : NOR2D1 port map( A1 => mult_239_n96, A2 => mult_239_n109, Z 
                           => m2_out_0_port);
   mult_239_U74 : INVD1 port map( A => m2_in_r_2_port, Z => mult_239_n106);
   mult_239_U73 : INVD1 port map( A => m2_in_r_0_port, Z => mult_239_n109);
   mult_239_U72 : INVD1 port map( A => mult_239_n1, Z => m2_out_14_port);
   mult_239_U71 : INVD1 port map( A => mult_239_n27, Z => mult_239_n108);
   mult_239_U70 : INVD1 port map( A => m2_in_r_5_port, Z => mult_239_n100);
   mult_239_U69 : INVD1 port map( A => m2_in_r_6_port, Z => mult_239_n98);
   mult_239_U68 : INVD1 port map( A => m2_in_r_4_port, Z => mult_239_n102);
   mult_239_U67 : INVD1 port map( A => m2_in_r_3_port, Z => mult_239_n104);
   mult_239_U66 : INVD1 port map( A => m2_in_r_1_port, Z => mult_239_n107);
   mult_239_U65 : INVD1 port map( A => mult_239_n15, Z => mult_239_n99);
   mult_239_U64 : INVD1 port map( A => mult_239_n17, Z => mult_239_n101);
   mult_239_U63 : INVD1 port map( A => mult_239_n19, Z => mult_239_n103);
   mult_239_U62 : INVD1 port map( A => mult_239_n21, Z => mult_239_n105);
   mult_239_U61 : INVD1 port map( A => m5_in_l_0, Z => mult_239_n96);
   mult_239_U22 : ADHALFDL port map( A => mult_239_n35, B => mult_239_n42, CO 
                           => mult_239_n28, S => mult_239_n29);
   mult_239_U20 : ADFULD1 port map( A => mult_239_n41, B => mult_239_n34, CI =>
                           mult_239_n27, CO => mult_239_n24, S => mult_239_n25)
                           ;
   mult_239_U19 : ADFULD1 port map( A => mult_239_n31, B => mult_239_n108, CI 
                           => mult_239_n33, CO => mult_239_n22, S => 
                           mult_239_n23);
   mult_239_U14 : ADHALFDL port map( A => mult_239_n47, B => mult_239_n40, CO 
                           => mult_239_n13, S => m2_out_1_port);
   mult_239_U13 : ADFULD1 port map( A => mult_239_n46, B => mult_239_n39, CI =>
                           mult_239_n13, CO => mult_239_n12, S => m2_out_2_port
                           );
   mult_239_U12 : ADFULD1 port map( A => mult_239_n45, B => mult_239_n38, CI =>
                           mult_239_n12, CO => mult_239_n11, S => m2_out_3_port
                           );
   mult_239_U11 : ADFULD1 port map( A => mult_239_n44, B => mult_239_n37, CI =>
                           mult_239_n11, CO => mult_239_n10, S => m2_out_4_port
                           );
   mult_239_U10 : ADFULD1 port map( A => mult_239_n43, B => mult_239_n36, CI =>
                           mult_239_n10, CO => mult_239_n9, S => m2_out_5_port)
                           ;
   mult_239_U9 : ADFULD1 port map( A => mult_239_n29, B => mult_239_n32, CI => 
                           mult_239_n9, CO => mult_239_n8, S => m2_out_6_port);
   mult_239_U8 : ADFULD1 port map( A => mult_239_n25, B => mult_239_n28, CI => 
                           mult_239_n8, CO => mult_239_n7, S => m2_out_7_port);
   mult_239_U7 : ADFULD1 port map( A => mult_239_n23, B => mult_239_n24, CI => 
                           mult_239_n7, CO => mult_239_n6, S => m2_out_8_port);
   mult_239_U6 : ADFULD1 port map( A => mult_239_n22, B => mult_239_n21, CI => 
                           mult_239_n6, CO => mult_239_n5, S => m2_out_9_port);
   mult_239_U5 : ADFULD1 port map( A => mult_239_n19, B => mult_239_n105, CI =>
                           mult_239_n5, CO => mult_239_n4, S => m2_out_10_port)
                           ;
   mult_239_U4 : ADFULD1 port map( A => mult_239_n17, B => mult_239_n103, CI =>
                           mult_239_n4, CO => mult_239_n3, S => m2_out_11_port)
                           ;
   mult_239_U3 : ADFULD1 port map( A => mult_239_n15, B => mult_239_n101, CI =>
                           mult_239_n3, CO => mult_239_n2, S => m2_out_12_port)
                           ;
   mult_239_U2 : ADFULD1 port map( A => mult_239_n30, B => mult_239_n99, CI => 
                           mult_239_n2, CO => mult_239_n1, S => m2_out_13_port)
                           ;

end flat_rtl_none_10;
