
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_TRA3 is

-- define attributes
attribute ENUM_ENCODING : STRING;

-- define any necessary types
type SIGNED is array (INTEGER range <>) of std_logic;

end CONV_PACK_TRA3;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture hier_rtl_none_10 of TRA3_DW_mult_tc_4 is

   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n29, n30, n31, n32, n33
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, product_0_port, product_1_port,
      product_2_port, product_3_port, product_4_port, product_5_port, 
      product_6_port, product_7_port, product_8_port, product_9_port, 
      product_10_port, product_11_port, product_12_port, n119, product_13_port,
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130 : std_logic;

begin
   product <= ( product_13_port, product_13_port, product_12_port, 
      product_11_port, product_10_port, product_9_port, product_8_port, 
      product_7_port, product_6_port, product_5_port, product_4_port, 
      product_3_port, product_2_port, product_1_port, product_0_port );
   
   U4 : ADFULD1 port map( A => n12, B => n46, CI => n3, CO => n2, S => 
                           product_12_port);
   U5 : ADFULD1 port map( A => n13, B => n14, CI => n4, CO => n3, S => 
                           product_11_port);
   U6 : ADFULD1 port map( A => n15, B => n18, CI => n5, CO => n4, S => 
                           product_10_port);
   U7 : ADFULD1 port map( A => n19, B => n24, CI => n6, CO => n5, S => 
                           product_9_port);
   U8 : ADFULD1 port map( A => n25, B => n30, CI => n7, CO => n6, S => 
                           product_8_port);
   U9 : ADFULD1 port map( A => n31, B => n36, CI => n8, CO => n7, S => 
                           product_7_port);
   U10 : ADFULD1 port map( A => n37, B => n40, CI => n9, CO => n8, S => 
                           product_6_port);
   U11 : ADFULD1 port map( A => n10, B => n43, CI => n41, CO => n9, S => 
                           product_5_port);
   U12 : ADFULD1 port map( A => n11, B => n58, CI => n45, CO => n10, S => 
                           product_4_port);
   U13 : ADHALFDL port map( A => n71, B => n66, CO => n11, S => product_3_port)
                           ;
   U14 : ADFULD1 port map( A => n51, B => n47, CI => n16, CO => n12, S => n13);
   U15 : ADFULD1 port map( A => n20, B => n48, CI => n17, CO => n14, S => n15);
   U16 : ADFULD1 port map( A => n52, B => n124, CI => n59, CO => n16, S => n17)
                           ;
   U17 : ADFULD1 port map( A => n26, B => n23, CI => n21, CO => n18, S => n19);
   U18 : ADFULD1 port map( A => n126, B => n60, CI => n53, CO => n20, S => n21)
                           ;
   U20 : ADFULD1 port map( A => n32, B => n29, CI => n27, CO => n24, S => n25);
   U21 : ADFULD1 port map( A => n128, B => n61, CI => n54, CO => n26, S => n27)
                           ;
   U23 : ADFULD1 port map( A => n38, B => n35, CI => n33, CO => n30, S => n31);
   U24 : ADFULD1 port map( A => n55, B => n62, CI => n67, CO => n32, S => n33);
   U26 : ADFULD1 port map( A => n42, B => n68, CI => n39, CO => n36, S => n37);
   U27 : ADFULD1 port map( A => n49, B => n56, CI => n63, CO => n38, S => n39);
   U28 : ADFULD1 port map( A => n64, B => n69, CI => n44, CO => n40, S => n41);
   U29 : ADHALFDL port map( A => n50, B => n57, CO => n42, S => n43);
   U30 : ADHALFDL port map( A => n65, B => n70, CO => n44, S => n45);
   U78 : INVD1 port map( A => a(3), Z => n119);
   U79 : INVD1 port map( A => n2, Z => product_13_port);
   U80 : INVD1 port map( A => b(4), Z => n123);
   U81 : INVD1 port map( A => b(3), Z => n125);
   U82 : INVD1 port map( A => b(2), Z => n127);
   U83 : INVD1 port map( A => n35, Z => n128);
   U84 : INVD1 port map( A => n29, Z => n126);
   U85 : INVD1 port map( A => n23, Z => n124);
   U86 : INVD1 port map( A => b(0), Z => n130);
   U87 : INVD1 port map( A => b(1), Z => n129);
   U88 : INVD1 port map( A => b(5), Z => n122);
   U89 : INVD1 port map( A => b(6), Z => n121);
   U90 : NOR2D1 port map( A1 => n119, A2 => n127, Z => product_2_port);
   U91 : NOR2D1 port map( A1 => n119, A2 => n129, Z => product_1_port);
   U92 : NOR2D1 port map( A1 => n119, A2 => n130, Z => product_0_port);
   U93 : NOR2D1 port map( A1 => n119, A2 => n125, Z => n71);
   U94 : NOR2D1 port map( A1 => n119, A2 => n123, Z => n70);
   U95 : NOR2D1 port map( A1 => n119, A2 => n122, Z => n69);
   U96 : NOR2D1 port map( A1 => n119, A2 => n121, Z => n68);
   U97 : NAN2D1 port map( A1 => b(7), A2 => a(0), Z => n67);
   U98 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n66);
   U99 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n65);
   U100 : NOR2D1 port map( A1 => n127, A2 => n119, Z => n64);
   U101 : NOR2D1 port map( A1 => n125, A2 => n119, Z => n63);
   U102 : NOR2D1 port map( A1 => n123, A2 => n119, Z => n62);
   U103 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n61);
   U104 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n60);
   U105 : NAN2D1 port map( A1 => a(3), A2 => b(7), Z => n59);
   U106 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n58);
   U107 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n57);
   U108 : NOR2D1 port map( A1 => n127, A2 => n119, Z => n56);
   U109 : NOR2D1 port map( A1 => n125, A2 => n119, Z => n55);
   U110 : NOR2D1 port map( A1 => n123, A2 => n119, Z => n54);
   U111 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n53);
   U112 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n52);
   U113 : NAN2D1 port map( A1 => a(4), A2 => b(7), Z => n51);
   U114 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n50);
   U115 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n49);
   U116 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n48);
   U117 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n47);
   U118 : NAN2D1 port map( A1 => a(5), A2 => b(7), Z => n46);
   U119 : NAN2D1 port map( A1 => a(5), A2 => b(2), Z => n35);
   U120 : NAN2D1 port map( A1 => a(5), A2 => b(3), Z => n29);
   U121 : NAN2D1 port map( A1 => a(5), A2 => b(4), Z => n23);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture hier_rtl_none_10 of TRA3_DW_mult_tc_3 is

   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n15, n17, n19
      , n21, n22, n23, n24, n25, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n96, n98, n99
      , n100, n101, n102, n103, n104, n105, n106, n107, n108, n109 : std_logic;

begin
   
   U2 : ADFULD1 port map( A => n30, B => n99, CI => n2, CO => n1, S => 
                           product(13));
   U3 : ADFULD1 port map( A => n15, B => n101, CI => n3, CO => n2, S => 
                           product(12));
   U4 : ADFULD1 port map( A => n17, B => n103, CI => n4, CO => n3, S => 
                           product(11));
   U5 : ADFULD1 port map( A => n19, B => n105, CI => n5, CO => n4, S => 
                           product(10));
   U6 : ADFULD1 port map( A => n22, B => n21, CI => n6, CO => n5, S => 
                           product(9));
   U7 : ADFULD1 port map( A => n23, B => n24, CI => n7, CO => n6, S => 
                           product(8));
   U8 : ADFULD1 port map( A => n25, B => n28, CI => n8, CO => n7, S => 
                           product(7));
   U9 : ADFULD1 port map( A => n29, B => n32, CI => n9, CO => n8, S => 
                           product(6));
   U10 : ADFULD1 port map( A => n43, B => n36, CI => n10, CO => n9, S => 
                           product(5));
   U11 : ADFULD1 port map( A => n44, B => n37, CI => n11, CO => n10, S => 
                           product(4));
   U12 : ADFULD1 port map( A => n45, B => n38, CI => n12, CO => n11, S => 
                           product(3));
   U13 : ADFULD1 port map( A => n46, B => n39, CI => n13, CO => n12, S => 
                           product(2));
   U14 : ADHALFDL port map( A => n47, B => n40, CO => n13, S => product(1));
   U19 : ADFULD1 port map( A => n31, B => n108, CI => n33, CO => n22, S => n23)
                           ;
   U20 : ADFULD1 port map( A => n41, B => n34, CI => n27, CO => n24, S => n25);
   U22 : ADHALFDL port map( A => n35, B => n42, CO => n28, S => n29);
   U61 : INVD1 port map( A => a(0), Z => n96);
   U62 : INVD1 port map( A => n21, Z => n105);
   U63 : INVD1 port map( A => n19, Z => n103);
   U64 : INVD1 port map( A => n17, Z => n101);
   U65 : INVD1 port map( A => n15, Z => n99);
   U66 : INVD1 port map( A => b(1), Z => n107);
   U67 : INVD1 port map( A => b(3), Z => n104);
   U68 : INVD1 port map( A => b(4), Z => n102);
   U69 : INVD1 port map( A => b(6), Z => n98);
   U70 : INVD1 port map( A => b(5), Z => n100);
   U71 : INVD1 port map( A => n27, Z => n108);
   U72 : INVD1 port map( A => n1, Z => product(14));
   U73 : INVD1 port map( A => b(0), Z => n109);
   U74 : INVD1 port map( A => b(2), Z => n106);
   U75 : NOR2D1 port map( A1 => n96, A2 => n109, Z => product(0));
   U76 : NOR2D1 port map( A1 => n96, A2 => n107, Z => n47);
   U77 : NOR2D1 port map( A1 => n96, A2 => n106, Z => n46);
   U78 : NOR2D1 port map( A1 => n96, A2 => n104, Z => n45);
   U79 : NOR2D1 port map( A1 => n96, A2 => n102, Z => n44);
   U80 : NOR2D1 port map( A1 => n96, A2 => n100, Z => n43);
   U81 : NOR2D1 port map( A1 => n96, A2 => n98, Z => n42);
   U82 : NAN2D1 port map( A1 => b(7), A2 => a(0), Z => n41);
   U83 : NOR2D1 port map( A1 => n109, A2 => n96, Z => n40);
   U84 : NOR2D1 port map( A1 => n107, A2 => n96, Z => n39);
   U85 : NOR2D1 port map( A1 => n106, A2 => n96, Z => n38);
   U86 : NOR2D1 port map( A1 => n104, A2 => n96, Z => n37);
   U87 : NOR2D1 port map( A1 => n102, A2 => n96, Z => n36);
   U88 : NOR2D1 port map( A1 => n100, A2 => n96, Z => n35);
   U89 : NOR2D1 port map( A1 => n98, A2 => n96, Z => n34);
   U90 : NAN2D1 port map( A1 => a(1), A2 => b(7), Z => n33);
   U91 : NOR2D1 port map( A1 => n109, A2 => n96, Z => n32);
   U92 : NOR2D1 port map( A1 => n106, A2 => n96, Z => n31);
   U93 : NAN2D1 port map( A1 => a(6), A2 => b(7), Z => n30);
   U94 : NAN2D1 port map( A1 => a(6), A2 => b(1), Z => n27);
   U95 : NAN2D1 port map( A1 => a(6), A2 => b(3), Z => n21);
   U96 : NAN2D1 port map( A1 => a(6), A2 => b(4), Z => n19);
   U97 : NAN2D1 port map( A1 => a(6), A2 => b(5), Z => n17);
   U98 : NAN2D1 port map( A1 => a(6), A2 => b(6), Z => n15);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture hier_rtl_none_10 of TRA3_DW_mult_tc_2 is

   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n20, n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107
      , n108, n109, n110, n111, n112, n113, n114, n115, n167, n168, n169, n170,
      n171, n172, n173, n174, n175, n176, n177, n178, n179 : std_logic;

begin
   
   U3 : ADFULD1 port map( A => n16, B => n17, CI => n3, CO => n2, S => 
                           product(13));
   U4 : ADFULD1 port map( A => n21, B => n18, CI => n4, CO => n3, S => 
                           product(12));
   U5 : ADFULD1 port map( A => n25, B => n22, CI => n5, CO => n4, S => 
                           product(11));
   U6 : ADFULD1 port map( A => n26, B => n29, CI => n6, CO => n5, S => 
                           product(10));
   U7 : ADFULD1 port map( A => n30, B => n35, CI => n7, CO => n6, S => 
                           product(9));
   U8 : ADFULD1 port map( A => n36, B => n43, CI => n8, CO => n7, S => 
                           product(8));
   U9 : ADFULD1 port map( A => n44, B => n51, CI => n9, CO => n8, S => 
                           product(7));
   U10 : ADFULD1 port map( A => n52, B => n57, CI => n10, CO => n9, S => 
                           product(6));
   U11 : ADFULD1 port map( A => n58, B => n61, CI => n11, CO => n10, S => 
                           product(5));
   U12 : ADFULD1 port map( A => n62, B => n65, CI => n12, CO => n11, S => 
                           product(4));
   U13 : ADFULD1 port map( A => n13, B => n68, CI => n66, CO => n12, S => 
                           product(3));
   U14 : ADFULD1 port map( A => n14, B => n100, CI => n70, CO => n13, S => 
                           product(2));
   U15 : ADHALFDL port map( A => n115, B => n108, CO => n14, S => product(1));
   U16 : ADFULD1 port map( A => n79, B => n168, CI => n72, CO => n15, S => n16)
                           ;
   U17 : ADFULD1 port map( A => n73, B => n170, CI => n20, CO => n17, S => n18)
                           ;
   U19 : ADFULD1 port map( A => n24, B => n74, CI => n27, CO => n21, S => n22);
   U21 : ADFULD1 port map( A => n28, B => n33, CI => n31, CO => n25, S => n26);
   U22 : ADFULD1 port map( A => n85, B => n80, CI => n75, CO => n27, S => n28);
   U23 : ADFULD1 port map( A => n37, B => n34, CI => n32, CO => n29, S => n30);
   U24 : ADFULD1 port map( A => n41, B => n93, CI => n39, CO => n31, S => n32);
   U25 : ADFULD1 port map( A => n81, B => n86, CI => n76, CO => n33, S => n34);
   U26 : ADFULD1 port map( A => n45, B => n40, CI => n38, CO => n35, S => n36);
   U27 : ADFULD1 port map( A => n42, B => n49, CI => n47, CO => n37, S => n38);
   U28 : ADFULD1 port map( A => n101, B => n87, CI => n77, CO => n39, S => n40)
                           ;
   U31 : ADFULD1 port map( A => n48, B => n53, CI => n46, CO => n43, S => n44);
   U32 : ADFULD1 port map( A => n55, B => n109, CI => n50, CO => n45, S => n46)
                           ;
   U33 : ADFULD1 port map( A => n83, B => n102, CI => n78, CO => n47, S => n48)
                           ;
   U34 : ADHALFDL port map( A => n95, B => n88, CO => n49, S => n50);
   U35 : ADFULD1 port map( A => n59, B => n56, CI => n54, CO => n51, S => n52);
   U36 : ADFULD1 port map( A => n96, B => n110, CI => n103, CO => n53, S => n54
                           );
   U37 : ADHALFDL port map( A => n84, B => n89, CO => n55, S => n56);
   U38 : ADFULD1 port map( A => n63, B => n111, CI => n60, CO => n57, S => n58)
                           ;
   U39 : ADFULD1 port map( A => n90, B => n97, CI => n104, CO => n59, S => n60)
                           ;
   U40 : ADFULD1 port map( A => n67, B => n112, CI => n64, CO => n61, S => n62)
                           ;
   U41 : ADFULD1 port map( A => n91, B => n98, CI => n105, CO => n63, S => n64)
                           ;
   U42 : ADFULD1 port map( A => n106, B => n113, CI => n69, CO => n65, S => n66
                           );
   U43 : ADHALFDL port map( A => n92, B => n99, CO => n67, S => n68);
   U44 : ADHALFDL port map( A => n107, B => n114, CO => n69, S => n70);
   U110 : INVD1 port map( A => a(0), Z => n167);
   U111 : INVD1 port map( A => b(2), Z => n174);
   U112 : INVD1 port map( A => b(1), Z => n175);
   U113 : INVD1 port map( A => b(3), Z => n173);
   U114 : INVD1 port map( A => b(0), Z => n176);
   U115 : INVD1 port map( A => b(4), Z => n172);
   U116 : INVD1 port map( A => b(6), Z => n169);
   U117 : INVD1 port map( A => b(5), Z => n171);
   U118 : INVD1 port map( A => n24, Z => n170);
   U119 : INVD1 port map( A => n20, Z => n168);
   U120 : EXOR3D1 port map( A1 => n2, A2 => n15, A3 => n177, Z => product(14));
   U121 : AND2D1 port map( A1 => a(7), A2 => b(7), Z => n177);
   U122 : NOR2D1 port map( A1 => n167, A2 => n176, Z => product(0));
   U123 : NOR2D1 port map( A1 => n167, A2 => n175, Z => n99);
   U124 : NOR2D1 port map( A1 => n167, A2 => n174, Z => n98);
   U125 : NOR2D1 port map( A1 => n167, A2 => n173, Z => n97);
   U126 : NOR2D1 port map( A1 => n167, A2 => n172, Z => n96);
   U127 : NOR2D1 port map( A1 => n167, A2 => n171, Z => n95);
   U128 : NAN2D1 port map( A1 => a(2), A2 => b(7), Z => n93);
   U129 : NOR2D1 port map( A1 => n176, A2 => n167, Z => n92);
   U130 : NOR2D1 port map( A1 => n175, A2 => n167, Z => n91);
   U131 : NOR2D1 port map( A1 => n174, A2 => n167, Z => n90);
   U132 : NOR2D1 port map( A1 => n173, A2 => n167, Z => n89);
   U133 : NOR2D1 port map( A1 => n172, A2 => n167, Z => n88);
   U134 : NOR2D1 port map( A1 => n171, A2 => n167, Z => n87);
   U135 : NOR2D1 port map( A1 => n167, A2 => n169, Z => n86);
   U136 : NAN2D1 port map( A1 => a(3), A2 => b(7), Z => n85);
   U137 : NOR2D1 port map( A1 => n176, A2 => n167, Z => n84);
   U138 : NOR2D1 port map( A1 => n175, A2 => n167, Z => n83);
   U139 : NOR2D1 port map( A1 => n173, A2 => n167, Z => n81);
   U140 : NOR2D1 port map( A1 => n172, A2 => n167, Z => n80);
   U141 : NAN2D1 port map( A1 => a(6), A2 => b(7), Z => n79);
   U142 : NAN2D1 port map( A1 => b(0), A2 => a(7), Z => n78);
   U143 : NAN2D1 port map( A1 => b(1), A2 => a(7), Z => n77);
   U144 : NAN2D1 port map( A1 => b(2), A2 => a(7), Z => n76);
   U145 : NAN2D1 port map( A1 => b(3), A2 => a(7), Z => n75);
   U146 : NAN2D1 port map( A1 => b(4), A2 => a(7), Z => n74);
   U147 : NAN2D1 port map( A1 => b(5), A2 => a(7), Z => n73);
   U148 : NAN2D1 port map( A1 => b(6), A2 => a(7), Z => n72);
   U149 : EXNOR2D1 port map( A1 => n178, A2 => n179, Z => n42);
   U150 : NAN2D1 port map( A1 => n179, A2 => n178, Z => n41);
   U151 : NAN2D1 port map( A1 => a(6), A2 => b(2), Z => n178);
   U152 : NAN2D1 port map( A1 => b(6), A2 => a(2), Z => n179);
   U153 : NAN2D1 port map( A1 => a(6), A2 => b(5), Z => n24);
   U154 : NAN2D1 port map( A1 => a(6), A2 => b(6), Z => n20);
   U155 : NOR2D1 port map( A1 => n167, A2 => n175, Z => n115);
   U156 : NOR2D1 port map( A1 => n167, A2 => n174, Z => n114);
   U157 : NOR2D1 port map( A1 => n167, A2 => n173, Z => n113);
   U158 : NOR2D1 port map( A1 => n167, A2 => n172, Z => n112);
   U159 : NOR2D1 port map( A1 => n167, A2 => n171, Z => n111);
   U160 : NOR2D1 port map( A1 => n167, A2 => n169, Z => n110);
   U161 : NAN2D1 port map( A1 => a(0), A2 => b(7), Z => n109);
   U162 : NOR2D1 port map( A1 => n176, A2 => n167, Z => n108);
   U163 : NOR2D1 port map( A1 => n175, A2 => n167, Z => n107);
   U164 : NOR2D1 port map( A1 => n174, A2 => n167, Z => n106);
   U165 : NOR2D1 port map( A1 => n173, A2 => n167, Z => n105);
   U166 : NOR2D1 port map( A1 => n172, A2 => n167, Z => n104);
   U167 : NOR2D1 port map( A1 => n171, A2 => n167, Z => n103);
   U168 : NOR2D1 port map( A1 => n169, A2 => n167, Z => n102);
   U169 : NAN2D1 port map( A1 => a(1), A2 => b(7), Z => n101);
   U170 : NOR2D1 port map( A1 => n176, A2 => n167, Z => n100);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture hier_rtl_none_10 of TRA3_DW_mult_tc_1 is

   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n28, n29, n30, n31, n32, n34, n35
      , n36, n37, n38, n39, n40, n41, n42, n43, n44, n46, n47, n48, n49, n50, 
      n51, n52, n53, n54, n55, n56, n57, n58, n59, n61, n62, n63, n64, n65, n67
      , n68, n69, n70, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130 : std_logic;

begin
   
   U3 : ADFULD1 port map( A => n14, B => n15, CI => n3, CO => n2, S => 
                           product(13));
   U4 : ADFULD1 port map( A => n17, B => n122, CI => n4, CO => n3, S => 
                           product(12));
   U5 : ADFULD1 port map( A => n18, B => n19, CI => n5, CO => n4, S => 
                           product(11));
   U6 : ADFULD1 port map( A => n20, B => n23, CI => n6, CO => n5, S => 
                           product(10));
   U7 : ADFULD1 port map( A => n24, B => n29, CI => n7, CO => n6, S => 
                           product(9));
   U8 : ADFULD1 port map( A => n30, B => n35, CI => n8, CO => n7, S => 
                           product(8));
   U9 : ADFULD1 port map( A => n36, B => n39, CI => n9, CO => n8, S => 
                           product(7));
   U10 : ADFULD1 port map( A => n40, B => n41, CI => n10, CO => n9, S => 
                           product(6));
   U11 : ADFULD1 port map( A => n42, B => n43, CI => n11, CO => n10, S => 
                           product(5));
   U12 : ADFULD1 port map( A => n12, B => n57, CI => n44, CO => n11, S => 
                           product(4));
   U13 : ADHALFDL port map( A => n70, B => n64, CO => n12, S => product(3));
   U16 : ADFULD1 port map( A => n46, B => n51, CI => n21, CO => n17, S => n18);
   U17 : ADFULD1 port map( A => n25, B => n58, CI => n22, CO => n19, S => n20);
   U18 : ADFULD1 port map( A => n52, B => n120, CI => n47, CO => n21, S => n22)
                           ;
   U19 : ADFULD1 port map( A => n31, B => n28, CI => n26, CO => n23, S => n24);
   U20 : ADFULD1 port map( A => n123, B => n53, CI => n48, CO => n25, S => n26)
                           ;
   U22 : ADFULD1 port map( A => n37, B => n34, CI => n32, CO => n29, S => n30);
   U23 : ADFULD1 port map( A => n65, B => n59, CI => n49, CO => n31, S => n32);
   U25 : ADFULD1 port map( A => n50, B => n54, CI => n38, CO => n35, S => n36);
   U28 : ADFULD1 port map( A => n55, B => n67, CI => n61, CO => n39, S => n40);
   U29 : ADFULD1 port map( A => n56, B => n68, CI => n62, CO => n41, S => n42);
   U30 : ADHALFDL port map( A => n63, B => n69, CO => n43, S => n44);
   U78 : INVD1 port map( A => a(3), Z => n119);
   U79 : INVD1 port map( A => n15, Z => n122);
   U80 : INVD1 port map( A => b(3), Z => n124);
   U81 : INVD1 port map( A => b(1), Z => n126);
   U82 : INVD1 port map( A => b(2), Z => n125);
   U83 : INVD1 port map( A => b(0), Z => n127);
   U84 : INVD1 port map( A => b(5), Z => n121);
   U85 : INVD1 port map( A => n34, Z => n123);
   U86 : INVD1 port map( A => n28, Z => n120);
   U87 : NOR2D1 port map( A1 => n119, A2 => n126, Z => product(2));
   U88 : NOR2D1 port map( A1 => n119, A2 => n127, Z => product(1));
   U89 : EXNOR3D1 port map( A1 => n2, A2 => n128, A3 => n14, Z => product(14));
   U90 : AND2D1 port map( A1 => a(7), A2 => b(7), Z => n128);
   U91 : NOR2D1 port map( A1 => n119, A2 => n125, Z => n70);
   U92 : NOR2D1 port map( A1 => n119, A2 => n124, Z => n69);
   U93 : NOR2M1D1 port map( A1 => b(4), A2 => n119, Z => n68);
   U94 : NOR2D1 port map( A1 => n119, A2 => n121, Z => n67);
   U95 : NAN2D1 port map( A1 => b(7), A2 => a(1), Z => n65);
   U96 : NOR2D1 port map( A1 => n127, A2 => n119, Z => n64);
   U97 : NOR2D1 port map( A1 => n126, A2 => n119, Z => n63);
   U98 : NOR2D1 port map( A1 => n125, A2 => n119, Z => n62);
   U99 : NOR2D1 port map( A1 => n124, A2 => n119, Z => n61);
   U100 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n59);
   U101 : NAN2D1 port map( A1 => a(3), A2 => b(7), Z => n58);
   U102 : NOR2D1 port map( A1 => n127, A2 => n119, Z => n57);
   U103 : NOR2D1 port map( A1 => n126, A2 => n119, Z => n56);
   U104 : NOR2D1 port map( A1 => n125, A2 => n119, Z => n55);
   U105 : NOR2D1 port map( A1 => n124, A2 => n119, Z => n54);
   U106 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n53);
   U107 : NOR2M1D1 port map( A1 => b(6), A2 => n119, Z => n52);
   U108 : NAN2D1 port map( A1 => a(4), A2 => b(7), Z => n51);
   U109 : NAN2D1 port map( A1 => a(7), A2 => b(0), Z => n50);
   U110 : NAN2D1 port map( A1 => a(7), A2 => b(1), Z => n49);
   U111 : NAN2D1 port map( A1 => b(2), A2 => a(7), Z => n48);
   U112 : NAN2D1 port map( A1 => b(3), A2 => a(7), Z => n47);
   U113 : NAN2D1 port map( A1 => b(4), A2 => a(7), Z => n46);
   U114 : EXNOR2D1 port map( A1 => n129, A2 => n130, Z => n38);
   U115 : NAN2D1 port map( A1 => n129, A2 => n130, Z => n37);
   U116 : NAN2D1 port map( A1 => b(6), A2 => a(1), Z => n130);
   U117 : NAN2D1 port map( A1 => a(3), A2 => b(4), Z => n129);
   U118 : NAN2D1 port map( A1 => a(4), A2 => b(4), Z => n34);
   U119 : NAN2D1 port map( A1 => a(3), A2 => b(6), Z => n28);
   U120 : NAN2D1 port map( A1 => b(5), A2 => a(7), Z => n15);
   U121 : AND2D1 port map( A1 => b(6), A2 => a(7), Z => n14);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture hier_rtl_none_10 of TRA3_DW_mult_tc_0 is

   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n23, n24, n25, n26, n27, n29, n30, n31, n32, n33
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, product_0_port, product_1_port,
      product_2_port, product_3_port, product_4_port, product_5_port, 
      product_6_port, product_7_port, product_8_port, product_9_port, 
      product_10_port, product_11_port, product_12_port, n119, product_13_port,
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130 : std_logic;

begin
   product <= ( product_13_port, product_13_port, product_12_port, 
      product_11_port, product_10_port, product_9_port, product_8_port, 
      product_7_port, product_6_port, product_5_port, product_4_port, 
      product_3_port, product_2_port, product_1_port, product_0_port );
   
   U4 : ADFULD1 port map( A => n12, B => n46, CI => n3, CO => n2, S => 
                           product_12_port);
   U5 : ADFULD1 port map( A => n13, B => n14, CI => n4, CO => n3, S => 
                           product_11_port);
   U6 : ADFULD1 port map( A => n15, B => n18, CI => n5, CO => n4, S => 
                           product_10_port);
   U7 : ADFULD1 port map( A => n19, B => n24, CI => n6, CO => n5, S => 
                           product_9_port);
   U8 : ADFULD1 port map( A => n25, B => n30, CI => n7, CO => n6, S => 
                           product_8_port);
   U9 : ADFULD1 port map( A => n31, B => n36, CI => n8, CO => n7, S => 
                           product_7_port);
   U10 : ADFULD1 port map( A => n37, B => n40, CI => n9, CO => n8, S => 
                           product_6_port);
   U11 : ADFULD1 port map( A => n10, B => n43, CI => n41, CO => n9, S => 
                           product_5_port);
   U12 : ADFULD1 port map( A => n11, B => n58, CI => n45, CO => n10, S => 
                           product_4_port);
   U13 : ADHALFDL port map( A => n71, B => n66, CO => n11, S => product_3_port)
                           ;
   U14 : ADFULD1 port map( A => n51, B => n47, CI => n16, CO => n12, S => n13);
   U15 : ADFULD1 port map( A => n20, B => n48, CI => n17, CO => n14, S => n15);
   U16 : ADFULD1 port map( A => n52, B => n124, CI => n59, CO => n16, S => n17)
                           ;
   U17 : ADFULD1 port map( A => n26, B => n23, CI => n21, CO => n18, S => n19);
   U18 : ADFULD1 port map( A => n126, B => n60, CI => n53, CO => n20, S => n21)
                           ;
   U20 : ADFULD1 port map( A => n32, B => n29, CI => n27, CO => n24, S => n25);
   U21 : ADFULD1 port map( A => n128, B => n61, CI => n54, CO => n26, S => n27)
                           ;
   U23 : ADFULD1 port map( A => n38, B => n35, CI => n33, CO => n30, S => n31);
   U24 : ADFULD1 port map( A => n55, B => n62, CI => n67, CO => n32, S => n33);
   U26 : ADFULD1 port map( A => n42, B => n68, CI => n39, CO => n36, S => n37);
   U27 : ADFULD1 port map( A => n49, B => n56, CI => n63, CO => n38, S => n39);
   U28 : ADFULD1 port map( A => n64, B => n69, CI => n44, CO => n40, S => n41);
   U29 : ADHALFDL port map( A => n50, B => n57, CO => n42, S => n43);
   U30 : ADHALFDL port map( A => n65, B => n70, CO => n44, S => n45);
   U78 : INVD1 port map( A => a(3), Z => n119);
   U79 : INVD1 port map( A => n2, Z => product_13_port);
   U80 : INVD1 port map( A => b(4), Z => n123);
   U81 : INVD1 port map( A => b(2), Z => n127);
   U82 : INVD1 port map( A => b(3), Z => n125);
   U83 : INVD1 port map( A => n35, Z => n128);
   U84 : INVD1 port map( A => n29, Z => n126);
   U85 : INVD1 port map( A => n23, Z => n124);
   U86 : INVD1 port map( A => b(1), Z => n129);
   U87 : INVD1 port map( A => b(0), Z => n130);
   U88 : INVD1 port map( A => b(5), Z => n122);
   U89 : INVD1 port map( A => b(6), Z => n121);
   U90 : NOR2D1 port map( A1 => n119, A2 => n127, Z => product_2_port);
   U91 : NOR2D1 port map( A1 => n119, A2 => n129, Z => product_1_port);
   U92 : NOR2D1 port map( A1 => n119, A2 => n130, Z => product_0_port);
   U93 : NOR2D1 port map( A1 => n119, A2 => n125, Z => n71);
   U94 : NOR2D1 port map( A1 => n119, A2 => n123, Z => n70);
   U95 : NOR2D1 port map( A1 => n119, A2 => n122, Z => n69);
   U96 : NOR2D1 port map( A1 => n119, A2 => n121, Z => n68);
   U97 : NAN2D1 port map( A1 => b(7), A2 => a(0), Z => n67);
   U98 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n66);
   U99 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n65);
   U100 : NOR2D1 port map( A1 => n127, A2 => n119, Z => n64);
   U101 : NOR2D1 port map( A1 => n125, A2 => n119, Z => n63);
   U102 : NOR2D1 port map( A1 => n123, A2 => n119, Z => n62);
   U103 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n61);
   U104 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n60);
   U105 : NAN2D1 port map( A1 => a(3), A2 => b(7), Z => n59);
   U106 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n58);
   U107 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n57);
   U108 : NOR2D1 port map( A1 => n127, A2 => n119, Z => n56);
   U109 : NOR2D1 port map( A1 => n125, A2 => n119, Z => n55);
   U110 : NOR2D1 port map( A1 => n123, A2 => n119, Z => n54);
   U111 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n53);
   U112 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n52);
   U113 : NAN2D1 port map( A1 => a(4), A2 => b(7), Z => n51);
   U114 : NOR2D1 port map( A1 => n130, A2 => n119, Z => n50);
   U115 : NOR2D1 port map( A1 => n129, A2 => n119, Z => n49);
   U116 : NOR2D1 port map( A1 => n122, A2 => n119, Z => n48);
   U117 : NOR2D1 port map( A1 => n121, A2 => n119, Z => n47);
   U118 : NAN2D1 port map( A1 => a(5), A2 => b(7), Z => n46);
   U119 : NAN2D1 port map( A1 => a(5), A2 => b(2), Z => n35);
   U120 : NAN2D1 port map( A1 => a(5), A2 => b(3), Z => n29);
   U121 : NAN2D1 port map( A1 => a(5), A2 => b(4), Z => n23);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture hier_rtl_none_10 of TRA3_DW01_add_3 is

   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, n1
      , n2, n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1_13 : ADFULD1 port map( A => A(13), B => B(13), CI => carry_13_port, CO =>
                           carry_14_port, S => SUM(13));
   U1_12 : ADFULD1 port map( A => A(12), B => B(12), CI => carry_12_port, CO =>
                           carry_13_port, S => SUM(12));
   U1_11 : ADFULD1 port map( A => A(11), B => B(11), CI => carry_11_port, CO =>
                           carry_12_port, S => SUM(11));
   U1_10 : ADFULD1 port map( A => A(10), B => B(10), CI => carry_10_port, CO =>
                           carry_11_port, S => SUM(10));
   U1_9 : ADFULD1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : ADFULD1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : ADFULD1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : ADFULD1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_14 : EXOR3D1 port map( A1 => A(14), A2 => B(14), A3 => carry_14_port, Z 
                           => SUM(14));
   U1 : OAI21M20D1 port map( A1 => n1, A2 => A(5), B => n2, Z => carry_6_port);
   U2 : OAI21D1 port map( A1 => A(5), A2 => n1, B => B(5), Z => n2);
   U3 : OAI21M20D1 port map( A1 => n3, A2 => A(4), B => n4, Z => n1);
   U4 : OAI21D1 port map( A1 => A(4), A2 => n3, B => B(4), Z => n4);
   U5 : OAI21M20D1 port map( A1 => n5, A2 => A(3), B => n6, Z => n3);
   U6 : OAI21D1 port map( A1 => A(3), A2 => n5, B => B(3), Z => n6);
   U7 : OAI21M20D1 port map( A1 => n7, A2 => A(2), B => n8, Z => n5);
   U8 : OAI21D1 port map( A1 => A(2), A2 => n7, B => B(2), Z => n8);
   U9 : OAI21M20D1 port map( A1 => A(1), A2 => B(1), B => n9, Z => n7);
   U10 : OAI211D1 port map( A1 => A(1), A2 => B(1), B => A(0), C => B(0), Z => 
                           n9);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture hier_rtl_none_10 of TRA3_DW01_add_1 is

   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_14_port, carry_13_port, carry_12_port, carry_11_port, 
      carry_10_port, carry_9_port, carry_8_port, carry_7_port, carry_6_port, n1
      , n2, n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1_13 : ADFULD1 port map( A => A(13), B => B(13), CI => carry_13_port, CO =>
                           carry_14_port, S => SUM(13));
   U1_12 : ADFULD1 port map( A => A(12), B => B(12), CI => carry_12_port, CO =>
                           carry_13_port, S => SUM(12));
   U1_11 : ADFULD1 port map( A => A(11), B => B(11), CI => carry_11_port, CO =>
                           carry_12_port, S => SUM(11));
   U1_10 : ADFULD1 port map( A => A(10), B => B(10), CI => carry_10_port, CO =>
                           carry_11_port, S => SUM(10));
   U1_9 : ADFULD1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : ADFULD1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : ADFULD1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : ADFULD1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_14 : EXOR3D1 port map( A1 => A(14), A2 => B(14), A3 => carry_14_port, Z 
                           => SUM(14));
   U1 : OAI21M20D1 port map( A1 => n1, A2 => A(5), B => n2, Z => carry_6_port);
   U2 : OAI21D1 port map( A1 => A(5), A2 => n1, B => B(5), Z => n2);
   U3 : OAI21M20D1 port map( A1 => n3, A2 => A(4), B => n4, Z => n1);
   U4 : OAI21D1 port map( A1 => A(4), A2 => n3, B => B(4), Z => n4);
   U5 : OAI21M20D1 port map( A1 => n5, A2 => A(3), B => n6, Z => n3);
   U6 : OAI21D1 port map( A1 => A(3), A2 => n5, B => B(3), Z => n6);
   U7 : OAI21M20D1 port map( A1 => n7, A2 => A(2), B => n8, Z => n5);
   U8 : OAI21D1 port map( A1 => A(2), A2 => n7, B => B(2), Z => n8);
   U9 : OAI21M20D1 port map( A1 => A(1), A2 => B(1), B => n9, Z => n7);
   U10 : OAI211D1 port map( A1 => A(1), A2 => B(1), B => A(0), C => B(0), Z => 
                           n9);

end hier_rtl_none_10;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_TRA3.all;

architecture hier_rtl_none_10 of TRA3 is

   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2D2
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVBD2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFERPQ1
      port( D, CEB, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component TRA3_DW_mult_tc_3
      port( a, b : in std_logic_vector (7 downto 0);  product : out 
            std_logic_vector (15 downto 0));
   end component;
   
   component TRA3_DW_mult_tc_2
      port( a, b : in std_logic_vector (7 downto 0);  product : out 
            std_logic_vector (15 downto 0));
   end component;
   
   component TRA3_DW_mult_tc_1
      port( a, b : in std_logic_vector (7 downto 0);  product : out 
            std_logic_vector (15 downto 0));
   end component;
   
   component TRA3_DW_mult_tc_0
      port( a : in std_logic_vector (6 downto 0);  b : in std_logic_vector (7 
            downto 0);  product : out std_logic_vector (14 downto 0));
   end component;
   
   component TRA3_DW_mult_tc_4
      port( a : in std_logic_vector (6 downto 0);  b : in std_logic_vector (7 
            downto 0);  product : out std_logic_vector (14 downto 0));
   end component;
   
   component TRA3_DW01_add_3
      port( A, B : in std_logic_vector (14 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (14 downto 0);  CO : out std_logic);
   end component;
   
   component TRA3_DW01_add_1
      port( A, B : in std_logic_vector (14 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (14 downto 0);  CO : out std_logic);
   end component;
   
   component OAI22M10D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal arx_i1_reg_7_port, arx_i1_reg_6_port, arx_i1_reg_5_port, 
      arx_i1_reg_4_port, arx_i1_reg_3_port, arx_i1_reg_2_port, 
      arx_i1_reg_1_port, arx_i1_reg_0_port, arx_r1_reg_14_port, 
      arx_r1_reg_13_port, arx_r1_reg_12_port, arx_r1_reg_11_port, 
      arx_r1_reg_10_port, arx_r1_reg_9_port, arx_r1_reg_8_port, 
      arx_r1_reg_7_port, arx_r1_reg_6_port, arx_r1_reg_5_port, 
      arx_r1_reg_4_port, arx_r1_reg_3_port, arx_r1_reg_2_port, 
      arx_r1_reg_1_port, arx_r1_reg_0_port, arx_r2_reg_14_port, 
      arx_r2_reg_13_port, arx_r2_reg_12_port, arx_r2_reg_11_port, 
      arx_r2_reg_10_port, arx_r2_reg_9_port, arx_r2_reg_8_port, 
      arx_r2_reg_7_port, arx_r2_reg_6_port, arx_r2_reg_5_port, 
      arx_r2_reg_4_port, arx_r2_reg_3_port, arx_r2_reg_2_port, 
      arx_r2_reg_1_port, arx_r2_reg_0_port, arx_r3_reg_14_port, 
      arx_r3_reg_13_port, arx_r3_reg_12_port, arx_r3_reg_11_port, 
      arx_r3_reg_10_port, arx_r3_reg_9_port, arx_r3_reg_8_port, 
      arx_r3_reg_7_port, arx_r3_reg_6_port, arx_r3_reg_5_port, 
      arx_r3_reg_4_port, arx_r3_reg_3_port, arx_r3_reg_2_port, 
      arx_r3_reg_1_port, arx_r3_reg_0_port, arx_r4_reg_14_port, 
      arx_r4_reg_13_port, arx_r4_reg_12_port, arx_r4_reg_11_port, 
      arx_r4_reg_10_port, arx_r4_reg_9_port, arx_r4_reg_8_port, 
      arx_r4_reg_7_port, arx_r4_reg_6_port, arx_r4_reg_5_port, 
      arx_r4_reg_4_port, arx_r4_reg_3_port, arx_r4_reg_2_port, 
      arx_r4_reg_1_port, arx_d1_reg_14_port, arx_d1_reg_13_port, 
      arx_d1_reg_12_port, arx_d1_reg_11_port, arx_d1_reg_10_port, 
      arx_d1_reg_9_port, arx_d1_reg_8_port, arx_d1_reg_7_port, 
      arx_d2_reg_14_port, arx_d2_reg_13_port, arx_d2_reg_12_port, 
      arx_d2_reg_11_port, arx_d2_reg_10_port, arx_d2_reg_9_port, 
      arx_d2_reg_8_port, arx_d2_reg_7_port, arx_state_reg_1_port, 
      arx_state_reg_0_port, m1_in_r_7_port, m1_in_r_6_port, m1_in_r_5_port, 
      m1_in_r_4_port, m1_in_r_3_port, m1_in_r_2_port, m1_in_r_1_port, 
      m1_in_r_0_port, m1_out_15, m1_out_13_port, m1_out_12_port, m1_out_11_port
      , m1_out_10_port, m1_out_9_port, m1_out_8_port, m1_out_7_port, 
      m1_out_6_port, m1_out_5_port, m1_out_4_port, m1_out_3_port, m1_out_2_port
      , m1_out_1_port, m1_out_0_port, m2_in_r_7_port, m2_in_r_6_port, 
      m2_in_r_5_port, m2_in_r_4_port, m2_in_r_3_port, m2_in_r_2_port, 
      m2_in_r_1_port, m2_in_r_0_port, m2_out_14_port, m2_out_13_port, 
      m2_out_12_port, m2_out_11_port, m2_out_10_port, m2_out_9_port, 
      m2_out_8_port, m2_out_7_port, m2_out_6_port, m2_out_5_port, m2_out_4_port
      , m2_out_3_port, m2_out_2_port, m2_out_1_port, m2_out_0_port, 
      m3_out_14_port, m3_out_13_port, m3_out_12_port, m3_out_11_port, 
      m3_out_10_port, m3_out_9_port, m3_out_8_port, m3_out_7_port, 
      m3_out_6_port, m3_out_5_port, m3_out_4_port, m3_out_3_port, m3_out_2_port
      , m3_out_1_port, m4_in_r_7_port, m4_in_r_6_port, m4_in_r_5_port, 
      m4_in_r_4_port, m4_in_r_3_port, m4_in_r_2_port, m4_in_r_1_port, 
      m4_in_r_0_port, m4_out_14_port, m4_out_13_port, m4_out_12_port, 
      m4_out_11_port, m4_out_10_port, m4_out_9_port, m4_out_8_port, 
      m4_out_7_port, m4_out_6_port, m4_out_5_port, m4_out_4_port, m4_out_3_port
      , m4_out_2_port, m4_out_1_port, m4_out_0_port, m5_in_l_0, m5_in_r_7_port,
      m5_in_r_6_port, m5_in_r_5_port, m5_in_r_4_port, m5_in_r_3_port, 
      m5_in_r_2_port, m5_in_r_1_port, m5_in_r_0_port, m5_out_15, m5_out_13_port
      , m5_out_12_port, m5_out_11_port, m5_out_10_port, m5_out_9_port, 
      m5_out_8_port, m5_out_7_port, m5_out_6_port, m5_out_5_port, m5_out_4_port
      , m5_out_3_port, m5_out_2_port, m5_out_1_port, m5_out_0_port, 
      a1_in_l_14_port, a1_in_l_13_port, a1_in_l_12_port, a1_in_l_11_port, 
      a1_in_l_10_port, a1_in_l_9_port, a1_in_l_8_port, a1_in_l_7_port, 
      a1_in_l_6_port, a1_in_l_5_port, a1_in_l_4_port, a1_in_l_3_port, 
      a1_in_l_2_port, a1_in_l_1_port, a1_in_l_0_port, a1_in_r_14_port, 
      a1_in_r_13_port, a1_in_r_12_port, a1_in_r_11_port, a1_in_r_10_port, 
      a1_in_r_9_port, a1_in_r_8_port, a1_in_r_7_port, a1_in_r_6_port, 
      a1_in_r_5_port, a1_in_r_4_port, a1_in_r_3_port, a1_in_r_2_port, 
      a1_in_r_1_port, a1_in_r_0_port, a1_out_7_port, a1_out_6_port, 
      a1_out_5_port, a1_out_4_port, a1_out_3_port, a1_out_2_port, a1_out_1_port
      , a1_out_0_port, a2_in_l_14_port, a2_in_l_13_port, a2_in_l_12_port, 
      a2_in_l_11_port, a2_in_l_10_port, a2_in_l_9_port, a2_in_l_8_port, 
      a2_in_l_7_port, a2_in_l_6_port, a2_in_l_5_port, a2_in_l_4_port, 
      a2_in_l_3_port, a2_in_l_2_port, a2_in_l_1_port, a2_in_l_0_port, 
      a2_in_r_14_port, a2_in_r_13_port, a2_in_r_12_port, a2_in_r_11_port, 
      a2_in_r_10_port, a2_in_r_9_port, a2_in_r_8_port, a2_in_r_7_port, 
      a2_in_r_6_port, a2_in_r_5_port, a2_in_r_4_port, a2_in_r_3_port, 
      a2_in_r_2_port, a2_in_r_1_port, a2_in_r_0_port, a2_out_7_port, 
      a2_out_6_port, a2_out_5_port, a2_out_4_port, a2_out_3_port, a2_out_2_port
      , a2_out_1_port, a2_out_0_port, state_0_port, N44, N45, N46, N47, N48, 
      N49, N50, N51, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115
      , N116, N117, N118, N119, N120, N121, N122, N123, net1801, n92, n94, n95,
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n1060, n1070, 
      n1080, n1090, n1100, n1110, n1120, n1130, n1140, n1150, n1160, n1170, 
      n1180, n1190, n1200, n1210, n1220, n1230, n124, n125, n126, n127, n129, 
      n130, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, 
      n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, 
      n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, 
      n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      add_416_C244_rn_carry_1_port, add_416_C244_rn_carry_2_port, 
      add_416_C244_rn_carry_3_port, add_416_C244_rn_carry_4_port, 
      add_416_C244_rn_carry_5_port, add_416_C244_rn_carry_6_port, 
      add_416_C244_rn_carry_7_port, add_416_C243_rn_carry_1_port, 
      add_416_C243_rn_carry_2_port, add_416_C243_rn_carry_3_port, 
      add_416_C243_rn_carry_4_port, add_416_C243_rn_carry_5_port, 
      add_416_C243_rn_carry_6_port, add_416_C243_rn_carry_7_port, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n_1037, 
      n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, 
      n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054 : 
      std_logic;

begin
   
   U149 : OAI21D1 port map( A1 => n193, A2 => n247, B => n92, Z => n132);
   U150 : AOI22D1 port map( A1 => n190, A2 => a1_out_7_port, B1 => 
                           m2_out_14_port, B2 => n177, Z => n92);
   U151 : OAI21D1 port map( A1 => n193, A2 => n246, B => n94, Z => n133);
   U152 : AOI22D1 port map( A1 => n190, A2 => a1_out_6_port, B1 => 
                           m2_out_13_port, B2 => n177, Z => n94);
   U153 : OAI21D1 port map( A1 => n193, A2 => n245, B => n95, Z => n134);
   U154 : AOI22D1 port map( A1 => n190, A2 => a1_out_5_port, B1 => 
                           m2_out_12_port, B2 => n177, Z => n95);
   U155 : OAI21D1 port map( A1 => n193, A2 => n244, B => n96, Z => n135);
   U156 : AOI22D1 port map( A1 => n190, A2 => a1_out_4_port, B1 => 
                           m2_out_11_port, B2 => n177, Z => n96);
   U157 : OAI21D1 port map( A1 => n193, A2 => n243, B => n97, Z => n136);
   U158 : AOI22D1 port map( A1 => n190, A2 => a1_out_3_port, B1 => 
                           m2_out_10_port, B2 => n177, Z => n97);
   U159 : OAI21D1 port map( A1 => n193, A2 => n242, B => n98, Z => n137);
   U160 : AOI22D1 port map( A1 => n189, A2 => a1_out_2_port, B1 => 
                           m2_out_9_port, B2 => n177, Z => n98);
   U161 : OAI21D1 port map( A1 => n193, A2 => n241, B => n99, Z => n138);
   U162 : AOI22D1 port map( A1 => n189, A2 => a1_out_1_port, B1 => 
                           m2_out_8_port, B2 => n177, Z => n99);
   U163 : OAI21D1 port map( A1 => n193, A2 => n240, B => n100, Z => n139);
   U164 : AOI22D1 port map( A1 => n189, A2 => a1_out_0_port, B1 => 
                           m2_out_7_port, B2 => n177, Z => n100);
   U165 : OAI21D1 port map( A1 => n193, A2 => n239, B => n102, Z => n147);
   U166 : AOI22D1 port map( A1 => a2_out_7_port, A2 => n189, B1 => 
                           m4_out_14_port, B2 => n177, Z => n102);
   U167 : OAI21D1 port map( A1 => n193, A2 => n238, B => n103, Z => n148);
   U168 : AOI22D1 port map( A1 => a2_out_6_port, A2 => n189, B1 => 
                           m4_out_13_port, B2 => n177, Z => n103);
   U169 : OAI21D1 port map( A1 => n193, A2 => n237, B => n104, Z => n149);
   U170 : AOI22D1 port map( A1 => a2_out_5_port, A2 => n189, B1 => 
                           m4_out_12_port, B2 => n177, Z => n104);
   U171 : OAI21D1 port map( A1 => n193, A2 => n236, B => n105, Z => n150);
   U172 : AOI22D1 port map( A1 => a2_out_4_port, A2 => n189, B1 => 
                           m4_out_11_port, B2 => n177, Z => n105);
   U173 : OAI21D1 port map( A1 => n193, A2 => n235, B => n1060, Z => n151);
   U174 : AOI22D1 port map( A1 => a2_out_3_port, A2 => n189, B1 => 
                           m4_out_10_port, B2 => n177, Z => n1060);
   U175 : OAI21D1 port map( A1 => n193, A2 => n234, B => n1070, Z => n152);
   U176 : AOI22D1 port map( A1 => a2_out_2_port, A2 => n189, B1 => 
                           m4_out_9_port, B2 => n177, Z => n1070);
   U177 : OAI21D1 port map( A1 => n193, A2 => n233, B => n1080, Z => n153);
   U178 : AOI22D1 port map( A1 => a2_out_1_port, A2 => n189, B1 => 
                           m4_out_8_port, B2 => n177, Z => n1080);
   U179 : OAI21D1 port map( A1 => n193, A2 => n232, B => n1090, Z => n154);
   U180 : AOI22D1 port map( A1 => a2_out_0_port, A2 => n189, B1 => 
                           m4_out_7_port, B2 => n177, Z => n1090);
   U181 : OAI21D1 port map( A1 => n193, A2 => n217, B => n1120, Z => n162);
   U182 : AOI22D1 port map( A1 => m1_out_0_port, A2 => n189, B1 => 
                           m5_out_0_port, B2 => n177, Z => n1120);
   U183 : OAI21D1 port map( A1 => n193, A2 => n216, B => n1130, Z => n163);
   U184 : AOI22D1 port map( A1 => m1_out_1_port, A2 => n189, B1 => 
                           m5_out_1_port, B2 => n177, Z => n1130);
   U185 : OAI21D1 port map( A1 => n193, A2 => n215, B => n1140, Z => n164);
   U186 : AOI22D1 port map( A1 => m1_out_2_port, A2 => n189, B1 => 
                           m5_out_2_port, B2 => n177, Z => n1140);
   U187 : OAI21D1 port map( A1 => n193, A2 => n214, B => n1150, Z => n165);
   U188 : AOI22D1 port map( A1 => m1_out_3_port, A2 => n189, B1 => 
                           m5_out_3_port, B2 => n177, Z => n1150);
   U189 : OAI21D1 port map( A1 => n193, A2 => n213, B => n1160, Z => n166);
   U190 : AOI22D1 port map( A1 => m1_out_4_port, A2 => n189, B1 => 
                           m5_out_4_port, B2 => n177, Z => n1160);
   U191 : OAI21D1 port map( A1 => n193, A2 => n212, B => n1170, Z => n167);
   U192 : AOI22D1 port map( A1 => m1_out_5_port, A2 => n189, B1 => 
                           m5_out_5_port, B2 => n177, Z => n1170);
   U193 : OAI21D1 port map( A1 => n193, A2 => n211, B => n1180, Z => n168);
   U194 : AOI22D1 port map( A1 => m1_out_6_port, A2 => n189, B1 => 
                           m5_out_6_port, B2 => n177, Z => n1180);
   U195 : OAI21D1 port map( A1 => n193, A2 => n210, B => n1190, Z => n169);
   U196 : AOI22D1 port map( A1 => m1_out_7_port, A2 => n189, B1 => 
                           m5_out_7_port, B2 => n177, Z => n1190);
   U197 : OAI21D1 port map( A1 => n193, A2 => n209, B => n1200, Z => n170);
   U198 : AOI22D1 port map( A1 => m1_out_8_port, A2 => n189, B1 => 
                           m5_out_8_port, B2 => n177, Z => n1200);
   U199 : OAI21D1 port map( A1 => n193, A2 => n208, B => n1210, Z => n171);
   U200 : AOI22D1 port map( A1 => m1_out_9_port, A2 => n189, B1 => 
                           m5_out_9_port, B2 => n177, Z => n1210);
   U201 : OAI21D1 port map( A1 => n193, A2 => n207, B => n1220, Z => n172);
   U202 : AOI22D1 port map( A1 => m1_out_10_port, A2 => n189, B1 => 
                           m5_out_10_port, B2 => n177, Z => n1220);
   U203 : OAI21D1 port map( A1 => n193, A2 => n206, B => n1230, Z => n173);
   U204 : AOI22D1 port map( A1 => m1_out_11_port, A2 => n189, B1 => 
                           m5_out_11_port, B2 => n177, Z => n1230);
   U205 : OAI21D1 port map( A1 => n193, A2 => n205, B => n124, Z => n174);
   U206 : AOI22D1 port map( A1 => m1_out_12_port, A2 => n190, B1 => 
                           m5_out_12_port, B2 => n177, Z => n124);
   U207 : OAI21D1 port map( A1 => n193, A2 => n204, B => n125, Z => n175);
   U208 : AOI22D1 port map( A1 => m1_out_13_port, A2 => n189, B1 => 
                           m5_out_13_port, B2 => n177, Z => n125);
   U209 : OAI21D1 port map( A1 => n193, A2 => n203, B => n126, Z => n176);
   U210 : AOI22D1 port map( A1 => m1_out_15, A2 => n189, B1 => m5_out_15, B2 =>
                           n177, Z => n126);
   U211 : OAI22M10D1 port map( A1 => arx_r4_reg_9_port, A2 => n1110, B1 => n234
                           , B2 => n179, Z => a2_in_r_9_port);
   U212 : OAI22M10D1 port map( A1 => arx_r4_reg_8_port, A2 => n188, B1 => n233,
                           B2 => n179, Z => a2_in_r_8_port);
   U213 : OAI22M10D1 port map( A1 => arx_r4_reg_7_port, A2 => n188, B1 => n232,
                           B2 => n179, Z => a2_in_r_7_port);
   U214 : OAI22M10D1 port map( A1 => arx_r4_reg_6_port, A2 => n188, B1 => n225,
                           B2 => n179, Z => a2_in_r_6_port);
   U215 : OAI22M10D1 port map( A1 => arx_r4_reg_5_port, A2 => n188, B1 => n226,
                           B2 => n179, Z => a2_in_r_5_port);
   U216 : OAI22M10D1 port map( A1 => arx_r4_reg_4_port, A2 => n188, B1 => n227,
                           B2 => n179, Z => a2_in_r_4_port);
   U217 : OAI22M10D1 port map( A1 => arx_r4_reg_3_port, A2 => n188, B1 => n228,
                           B2 => n179, Z => a2_in_r_3_port);
   U218 : OAI22M10D1 port map( A1 => arx_r4_reg_2_port, A2 => n188, B1 => n229,
                           B2 => n179, Z => a2_in_r_2_port);
   U219 : OAI22M10D1 port map( A1 => arx_r4_reg_1_port, A2 => n188, B1 => n230,
                           B2 => n179, Z => a2_in_r_1_port);
   U220 : OAI22M10D1 port map( A1 => arx_r4_reg_14_port, A2 => n188, B1 => n239
                           , B2 => n179, Z => a2_in_r_14_port);
   U221 : OAI22M10D1 port map( A1 => arx_r4_reg_13_port, A2 => n1110, B1 => 
                           n238, B2 => n179, Z => a2_in_r_13_port);
   U222 : OAI22M10D1 port map( A1 => arx_r4_reg_12_port, A2 => n1110, B1 => 
                           n237, B2 => n179, Z => a2_in_r_12_port);
   U223 : OAI22M10D1 port map( A1 => arx_r4_reg_11_port, A2 => n1110, B1 => 
                           n236, B2 => n179, Z => a2_in_r_11_port);
   U224 : OAI22M10D1 port map( A1 => arx_r4_reg_10_port, A2 => n1110, B1 => 
                           n235, B2 => n179, Z => a2_in_r_10_port);
   U226 : OAI22D1 port map( A1 => n188, A2 => n234, B1 => n242, B2 => n179, Z 
                           => a1_in_r_9_port);
   U227 : OAI22D1 port map( A1 => n188, A2 => n233, B1 => n241, B2 => n179, Z 
                           => a1_in_r_8_port);
   U228 : OAI22D1 port map( A1 => n188, A2 => n232, B1 => n240, B2 => n179, Z 
                           => a1_in_r_7_port);
   U229 : OAI22D1 port map( A1 => n188, A2 => n225, B1 => n218, B2 => n179, Z 
                           => a1_in_r_6_port);
   U230 : OAI22D1 port map( A1 => n188, A2 => n226, B1 => n219, B2 => n179, Z 
                           => a1_in_r_5_port);
   U231 : OAI22D1 port map( A1 => n188, A2 => n227, B1 => n220, B2 => n179, Z 
                           => a1_in_r_4_port);
   U232 : OAI22D1 port map( A1 => n188, A2 => n228, B1 => n221, B2 => n179, Z 
                           => a1_in_r_3_port);
   U233 : OAI22D1 port map( A1 => n188, A2 => n229, B1 => n222, B2 => n179, Z 
                           => a1_in_r_2_port);
   U234 : OAI22D1 port map( A1 => n188, A2 => n230, B1 => n223, B2 => n179, Z 
                           => a1_in_r_1_port);
   U235 : OAI22D1 port map( A1 => n1110, A2 => n239, B1 => n247, B2 => n179, Z 
                           => a1_in_r_14_port);
   U236 : OAI22D1 port map( A1 => n1110, A2 => n238, B1 => n246, B2 => n179, Z 
                           => a1_in_r_13_port);
   U237 : OAI22D1 port map( A1 => n1110, A2 => n237, B1 => n245, B2 => n179, Z 
                           => a1_in_r_12_port);
   U238 : OAI22D1 port map( A1 => n1110, A2 => n236, B1 => n244, B2 => n179, Z 
                           => a1_in_r_11_port);
   U239 : OAI22D1 port map( A1 => n1110, A2 => n235, B1 => n243, B2 => n179, Z 
                           => a1_in_r_10_port);
   U240 : OAI22D1 port map( A1 => n188, A2 => n231, B1 => n224, B2 => n179, Z 
                           => a1_in_r_0_port);
   U241 : OAI22M10D1 port map( A1 => arx_i1_reg_2_port, A2 => n179, B1 => n1110
                           , B2 => n242, Z => a1_in_l_9_port);
   U242 : OAI22M10D1 port map( A1 => arx_i1_reg_1_port, A2 => n179, B1 => n1110
                           , B2 => n241, Z => a1_in_l_8_port);
   U243 : OAI22M10D1 port map( A1 => arx_i1_reg_0_port, A2 => n179, B1 => n188,
                           B2 => n240, Z => a1_in_l_7_port);
   U244 : OAI22M10D1 port map( A1 => arx_i1_reg_7_port, A2 => n179, B1 => n1110
                           , B2 => n247, Z => a1_in_l_14_port);
   U245 : OAI22M10D1 port map( A1 => arx_i1_reg_6_port, A2 => n179, B1 => n1110
                           , B2 => n246, Z => a1_in_l_13_port);
   U246 : OAI22M10D1 port map( A1 => arx_i1_reg_5_port, A2 => n179, B1 => n1110
                           , B2 => n245, Z => a1_in_l_12_port);
   U247 : OAI22M10D1 port map( A1 => arx_i1_reg_4_port, A2 => n179, B1 => n1110
                           , B2 => n244, Z => a1_in_l_11_port);
   U248 : OAI22M10D1 port map( A1 => arx_i1_reg_3_port, A2 => n179, B1 => n1110
                           , B2 => n243, Z => a1_in_l_10_port);
   add_244 : TRA3_DW01_add_1 port map( A(14) => a2_in_l_14_port, A(13) => 
                           a2_in_l_13_port, A(12) => a2_in_l_12_port, A(11) => 
                           a2_in_l_11_port, A(10) => a2_in_l_10_port, A(9) => 
                           a2_in_l_9_port, A(8) => a2_in_l_8_port, A(7) => 
                           a2_in_l_7_port, A(6) => a2_in_l_6_port, A(5) => 
                           a2_in_l_5_port, A(4) => a2_in_l_4_port, A(3) => 
                           a2_in_l_3_port, A(2) => a2_in_l_2_port, A(1) => 
                           a2_in_l_1_port, A(0) => a2_in_l_0_port, B(14) => 
                           a2_in_r_14_port, B(13) => a2_in_r_13_port, B(12) => 
                           a2_in_r_12_port, B(11) => a2_in_r_11_port, B(10) => 
                           a2_in_r_10_port, B(9) => a2_in_r_9_port, B(8) => 
                           a2_in_r_8_port, B(7) => a2_in_r_7_port, B(6) => 
                           a2_in_r_6_port, B(5) => a2_in_r_5_port, B(4) => 
                           a2_in_r_4_port, B(3) => a2_in_r_3_port, B(2) => 
                           a2_in_r_2_port, B(1) => a2_in_r_1_port, B(0) => 
                           a2_in_r_0_port, CI => net1801, SUM(14) => N123, 
                           SUM(13) => N122, SUM(12) => N121, SUM(11) => N120, 
                           SUM(10) => N119, SUM(9) => N118, SUM(8) => N117, 
                           SUM(7) => N116, SUM(6) => N115, SUM(5) => n_1037, 
                           SUM(4) => n_1038, SUM(3) => n_1039, SUM(2) => n_1040
                           , SUM(1) => n_1041, SUM(0) => n_1042, CO => n_1043);
   add_243 : TRA3_DW01_add_3 port map( A(14) => a1_in_l_14_port, A(13) => 
                           a1_in_l_13_port, A(12) => a1_in_l_12_port, A(11) => 
                           a1_in_l_11_port, A(10) => a1_in_l_10_port, A(9) => 
                           a1_in_l_9_port, A(8) => a1_in_l_8_port, A(7) => 
                           a1_in_l_7_port, A(6) => a1_in_l_6_port, A(5) => 
                           a1_in_l_5_port, A(4) => a1_in_l_4_port, A(3) => 
                           a1_in_l_3_port, A(2) => a1_in_l_2_port, A(1) => 
                           a1_in_l_1_port, A(0) => a1_in_l_0_port, B(14) => 
                           a1_in_r_14_port, B(13) => a1_in_r_13_port, B(12) => 
                           a1_in_r_12_port, B(11) => a1_in_r_11_port, B(10) => 
                           a1_in_r_10_port, B(9) => a1_in_r_9_port, B(8) => 
                           a1_in_r_8_port, B(7) => a1_in_r_7_port, B(6) => 
                           a1_in_r_6_port, B(5) => a1_in_r_5_port, B(4) => 
                           a1_in_r_4_port, B(3) => a1_in_r_3_port, B(2) => 
                           a1_in_r_2_port, B(1) => a1_in_r_1_port, B(0) => 
                           a1_in_r_0_port, CI => net1801, SUM(14) => N114, 
                           SUM(13) => N113, SUM(12) => N112, SUM(11) => N111, 
                           SUM(10) => N110, SUM(9) => N109, SUM(8) => N108, 
                           SUM(7) => N107, SUM(6) => N106, SUM(5) => n_1044, 
                           SUM(4) => n_1045, SUM(3) => n_1046, SUM(2) => n_1047
                           , SUM(1) => n_1048, SUM(0) => n_1049, CO => n_1050);
   mult_238 : TRA3_DW_mult_tc_4 port map( a(6) => net1801, a(5) => n193, a(4) 
                           => n193, a(3) => n193, a(2) => net1801, a(1) => 
                           net1801, a(0) => n193, b(7) => m1_in_r_7_port, b(6) 
                           => m1_in_r_6_port, b(5) => m1_in_r_5_port, b(4) => 
                           m1_in_r_4_port, b(3) => m1_in_r_3_port, b(2) => 
                           m1_in_r_2_port, b(1) => m1_in_r_1_port, b(0) => 
                           m1_in_r_0_port, product(14) => m1_out_15, 
                           product(13) => m1_out_13_port, product(12) => 
                           m1_out_12_port, product(11) => m1_out_11_port, 
                           product(10) => m1_out_10_port, product(9) => 
                           m1_out_9_port, product(8) => m1_out_8_port, 
                           product(7) => m1_out_7_port, product(6) => 
                           m1_out_6_port, product(5) => m1_out_5_port, 
                           product(4) => m1_out_4_port, product(3) => 
                           m1_out_3_port, product(2) => m1_out_2_port, 
                           product(1) => m1_out_1_port, product(0) => 
                           m1_out_0_port);
   mult_242 : TRA3_DW_mult_tc_0 port map( a(6) => net1801, a(5) => m5_in_l_0, 
                           a(4) => m5_in_l_0, a(3) => m5_in_l_0, a(2) => 
                           net1801, a(1) => net1801, a(0) => m5_in_l_0, b(7) =>
                           m5_in_r_7_port, b(6) => m5_in_r_6_port, b(5) => 
                           m5_in_r_5_port, b(4) => m5_in_r_4_port, b(3) => 
                           m5_in_r_3_port, b(2) => m5_in_r_2_port, b(1) => 
                           m5_in_r_1_port, b(0) => m5_in_r_0_port, product(14) 
                           => m5_out_15, product(13) => m5_out_13_port, 
                           product(12) => m5_out_12_port, product(11) => 
                           m5_out_11_port, product(10) => m5_out_10_port, 
                           product(9) => m5_out_9_port, product(8) => 
                           m5_out_8_port, product(7) => m5_out_7_port, 
                           product(6) => m5_out_6_port, product(5) => 
                           m5_out_5_port, product(4) => m5_out_4_port, 
                           product(3) => m5_out_3_port, product(2) => 
                           m5_out_2_port, product(1) => m5_out_1_port, 
                           product(0) => m5_out_0_port);
   mult_240 : TRA3_DW_mult_tc_1 port map( a(7) => m5_in_l_0, a(6) => net1801, 
                           a(5) => net1801, a(4) => m5_in_l_0, a(3) => 
                           m5_in_l_0, a(2) => net1801, a(1) => m5_in_l_0, a(0) 
                           => net1801, b(7) => m4_in_r_7_port, b(6) => 
                           m4_in_r_6_port, b(5) => m4_in_r_5_port, b(4) => 
                           m4_in_r_4_port, b(3) => m4_in_r_3_port, b(2) => 
                           m4_in_r_2_port, b(1) => m4_in_r_1_port, b(0) => 
                           m4_in_r_0_port, product(15) => n_1051, product(14) 
                           => m3_out_14_port, product(13) => m3_out_13_port, 
                           product(12) => m3_out_12_port, product(11) => 
                           m3_out_11_port, product(10) => m3_out_10_port, 
                           product(9) => m3_out_9_port, product(8) => 
                           m3_out_8_port, product(7) => m3_out_7_port, 
                           product(6) => m3_out_6_port, product(5) => 
                           m3_out_5_port, product(4) => m3_out_4_port, 
                           product(3) => m3_out_3_port, product(2) => 
                           m3_out_2_port, product(1) => m3_out_1_port, 
                           product(0) => n_1052);
   mult_241 : TRA3_DW_mult_tc_2 port map( a(7) => m5_in_l_0, a(6) => m5_in_l_0,
                           a(5) => net1801, a(4) => net1801, a(3) => m5_in_l_0,
                           a(2) => m5_in_l_0, a(1) => m5_in_l_0, a(0) => 
                           m5_in_l_0, b(7) => m4_in_r_7_port, b(6) => 
                           m4_in_r_6_port, b(5) => m4_in_r_5_port, b(4) => 
                           m4_in_r_4_port, b(3) => m4_in_r_3_port, b(2) => 
                           m4_in_r_2_port, b(1) => m4_in_r_1_port, b(0) => 
                           m4_in_r_0_port, product(15) => n_1053, product(14) 
                           => m4_out_14_port, product(13) => m4_out_13_port, 
                           product(12) => m4_out_12_port, product(11) => 
                           m4_out_11_port, product(10) => m4_out_10_port, 
                           product(9) => m4_out_9_port, product(8) => 
                           m4_out_8_port, product(7) => m4_out_7_port, 
                           product(6) => m4_out_6_port, product(5) => 
                           m4_out_5_port, product(4) => m4_out_4_port, 
                           product(3) => m4_out_3_port, product(2) => 
                           m4_out_2_port, product(1) => m4_out_1_port, 
                           product(0) => m4_out_0_port);
   mult_239 : TRA3_DW_mult_tc_3 port map( a(7) => net1801, a(6) => m5_in_l_0, 
                           a(5) => net1801, a(4) => net1801, a(3) => net1801, 
                           a(2) => net1801, a(1) => m5_in_l_0, a(0) => 
                           m5_in_l_0, b(7) => m2_in_r_7_port, b(6) => 
                           m2_in_r_6_port, b(5) => m2_in_r_5_port, b(4) => 
                           m2_in_r_4_port, b(3) => m2_in_r_3_port, b(2) => 
                           m2_in_r_2_port, b(1) => m2_in_r_1_port, b(0) => 
                           m2_in_r_0_port, product(15) => n_1054, product(14) 
                           => m2_out_14_port, product(13) => m2_out_13_port, 
                           product(12) => m2_out_12_port, product(11) => 
                           m2_out_11_port, product(10) => m2_out_10_port, 
                           product(9) => m2_out_9_port, product(8) => 
                           m2_out_8_port, product(7) => m2_out_7_port, 
                           product(6) => m2_out_6_port, product(5) => 
                           m2_out_5_port, product(4) => m2_out_4_port, 
                           product(3) => m2_out_3_port, product(2) => 
                           m2_out_2_port, product(1) => m2_out_1_port, 
                           product(0) => m2_out_0_port);
   arx_r1_reg_reg_14_inst : DFFRPQ1 port map( D => n176, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_14_port);
   arx_r4_reg_reg_14_inst : DFERPQ1 port map( D => m3_out_14_port, CEB => n1100
                           , CK => clock, RB => resetn, Q => arx_r4_reg_14_port
                           );
   arx_i1_reg_reg_7_inst : DFERPQ1 port map( D => data_in(7), CEB => n127, CK 
                           => clock, RB => resetn, Q => arx_i1_reg_7_port);
   arx_r2_reg_reg_14_inst : DFFRPQ1 port map( D => n132, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_14_port);
   arx_r3_reg_reg_14_inst : DFFRPQ1 port map( D => n147, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_14_port);
   arx_r1_reg_reg_13_inst : DFFRPQ1 port map( D => n175, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_13_port);
   arx_r4_reg_reg_13_inst : DFERPQ1 port map( D => m3_out_13_port, CEB => n1100
                           , CK => clock, RB => resetn, Q => arx_r4_reg_13_port
                           );
   arx_i1_reg_reg_6_inst : DFERPQ1 port map( D => data_in(6), CEB => n127, CK 
                           => clock, RB => resetn, Q => arx_i1_reg_6_port);
   arx_r2_reg_reg_13_inst : DFFRPQ1 port map( D => n133, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_13_port);
   arx_r3_reg_reg_13_inst : DFFRPQ1 port map( D => n148, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_13_port);
   arx_r1_reg_reg_12_inst : DFFRPQ1 port map( D => n174, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_12_port);
   arx_r4_reg_reg_12_inst : DFERPQ1 port map( D => m3_out_12_port, CEB => n1100
                           , CK => clock, RB => resetn, Q => arx_r4_reg_12_port
                           );
   arx_i1_reg_reg_5_inst : DFERPQ1 port map( D => data_in(5), CEB => n127, CK 
                           => clock, RB => resetn, Q => arx_i1_reg_5_port);
   arx_r2_reg_reg_12_inst : DFFRPQ1 port map( D => n134, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_12_port);
   arx_r3_reg_reg_12_inst : DFFRPQ1 port map( D => n149, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_12_port);
   arx_r1_reg_reg_11_inst : DFFRPQ1 port map( D => n173, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_11_port);
   arx_r4_reg_reg_11_inst : DFERPQ1 port map( D => m3_out_11_port, CEB => n1100
                           , CK => clock, RB => resetn, Q => arx_r4_reg_11_port
                           );
   arx_i1_reg_reg_4_inst : DFERPQ1 port map( D => data_in(4), CEB => n127, CK 
                           => clock, RB => resetn, Q => arx_i1_reg_4_port);
   arx_r2_reg_reg_11_inst : DFFRPQ1 port map( D => n135, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_11_port);
   arx_r3_reg_reg_11_inst : DFFRPQ1 port map( D => n150, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_11_port);
   arx_r1_reg_reg_10_inst : DFFRPQ1 port map( D => n172, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_10_port);
   arx_r4_reg_reg_10_inst : DFERPQ1 port map( D => m3_out_10_port, CEB => n1100
                           , CK => clock, RB => resetn, Q => arx_r4_reg_10_port
                           );
   arx_i1_reg_reg_3_inst : DFERPQ1 port map( D => data_in(3), CEB => n127, CK 
                           => clock, RB => resetn, Q => arx_i1_reg_3_port);
   arx_r2_reg_reg_10_inst : DFFRPQ1 port map( D => n136, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_10_port);
   arx_r3_reg_reg_10_inst : DFFRPQ1 port map( D => n151, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_10_port);
   arx_r1_reg_reg_9_inst : DFFRPQ1 port map( D => n171, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_9_port);
   arx_r4_reg_reg_9_inst : DFERPQ1 port map( D => m3_out_9_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_9_port);
   arx_i1_reg_reg_2_inst : DFERPQ1 port map( D => data_in(2), CEB => n127, CK 
                           => clock, RB => resetn, Q => arx_i1_reg_2_port);
   arx_r2_reg_reg_9_inst : DFFRPQ1 port map( D => n137, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_9_port);
   arx_r3_reg_reg_9_inst : DFFRPQ1 port map( D => n152, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_9_port);
   arx_r1_reg_reg_8_inst : DFFRPQ1 port map( D => n170, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_8_port);
   arx_r4_reg_reg_8_inst : DFERPQ1 port map( D => m3_out_8_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_8_port);
   arx_i1_reg_reg_1_inst : DFERPQ1 port map( D => data_in(1), CEB => n127, CK 
                           => clock, RB => resetn, Q => arx_i1_reg_1_port);
   arx_r2_reg_reg_8_inst : DFFRPQ1 port map( D => n138, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_8_port);
   arx_r3_reg_reg_8_inst : DFFRPQ1 port map( D => n153, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_8_port);
   arx_r1_reg_reg_7_inst : DFFRPQ1 port map( D => n169, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_7_port);
   arx_r4_reg_reg_7_inst : DFERPQ1 port map( D => m3_out_7_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_7_port);
   arx_i1_reg_reg_0_inst : DFERPQ1 port map( D => data_in(0), CEB => n127, CK 
                           => clock, RB => resetn, Q => arx_i1_reg_0_port);
   arx_r2_reg_reg_7_inst : DFFRPQ1 port map( D => n139, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_7_port);
   arx_r3_reg_reg_7_inst : DFFRPQ1 port map( D => n154, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_7_port);
   arx_d1_reg_reg_14_inst : DFERPQ1 port map( D => a1_out_7_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d1_reg_14_port);
   arx_d3_reg_reg_14_inst : DFERPQ1 port map( D => arx_d2_reg_14_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => N51);
   arx_d3_reg_reg_13_inst : DFERPQ1 port map( D => arx_d2_reg_13_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => N50);
   arx_d1_reg_reg_13_inst : DFERPQ1 port map( D => a1_out_6_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d1_reg_13_port);
   arx_r1_reg_reg_6_inst : DFFRPQ1 port map( D => n168, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_6_port);
   arx_r4_reg_reg_6_inst : DFERPQ1 port map( D => m3_out_6_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_6_port);
   arx_r2_reg_reg_6_inst : DFFRPQ1 port map( D => n140, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_6_port);
   arx_d1_reg_reg_12_inst : DFERPQ1 port map( D => a1_out_5_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d1_reg_12_port);
   arx_r3_reg_reg_6_inst : DFFRPQ1 port map( D => n155, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_6_port);
   arx_r4_reg_reg_5_inst : DFERPQ1 port map( D => m3_out_5_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_5_port);
   arx_r1_reg_reg_5_inst : DFFRPQ1 port map( D => n167, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_5_port);
   arx_d3_reg_reg_12_inst : DFERPQ1 port map( D => arx_d2_reg_12_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => N49);
   arx_r2_reg_reg_5_inst : DFFRPQ1 port map( D => n141, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_5_port);
   arx_r3_reg_reg_5_inst : DFFRPQ1 port map( D => n156, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_5_port);
   arx_d3_reg_reg_9_inst : DFERPQ1 port map( D => arx_d2_reg_9_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => N46);
   arx_d1_reg_reg_11_inst : DFERPQ1 port map( D => a1_out_4_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d1_reg_11_port);
   arx_d3_reg_reg_8_inst : DFERPQ1 port map( D => arx_d2_reg_8_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => N45);
   arx_d3_reg_reg_10_inst : DFERPQ1 port map( D => arx_d2_reg_10_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => N47);
   arx_d3_reg_reg_11_inst : DFERPQ1 port map( D => arx_d2_reg_11_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => N48);
   arx_d3_reg_reg_7_inst : DFERPQ1 port map( D => arx_d2_reg_7_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => N44);
   arx_r4_reg_reg_4_inst : DFERPQ1 port map( D => m3_out_4_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_4_port);
   arx_r1_reg_reg_4_inst : DFFRPQ1 port map( D => n166, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_4_port);
   arx_d1_reg_reg_10_inst : DFERPQ1 port map( D => a1_out_3_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d1_reg_10_port);
   arx_r2_reg_reg_4_inst : DFFRPQ1 port map( D => n142, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_4_port);
   arx_r3_reg_reg_4_inst : DFFRPQ1 port map( D => n157, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_4_port);
   arx_r4_reg_reg_3_inst : DFERPQ1 port map( D => m3_out_3_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_3_port);
   arx_r1_reg_reg_3_inst : DFFRPQ1 port map( D => n165, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_3_port);
   arx_r2_reg_reg_3_inst : DFFRPQ1 port map( D => n143, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_3_port);
   arx_r3_reg_reg_3_inst : DFFRPQ1 port map( D => n158, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_3_port);
   arx_d2_reg_reg_14_inst : DFERPQ1 port map( D => arx_d1_reg_14_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => 
                           arx_d2_reg_14_port);
   arx_d1_reg_reg_9_inst : DFERPQ1 port map( D => a1_out_2_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d1_reg_9_port);
   arx_d1_reg_reg_8_inst : DFERPQ1 port map( D => a1_out_1_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d1_reg_8_port);
   arx_d1_reg_reg_7_inst : DFERPQ1 port map( D => a1_out_0_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => arx_d1_reg_7_port);
   arx_r4_reg_reg_2_inst : DFERPQ1 port map( D => m3_out_2_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_2_port);
   arx_r1_reg_reg_2_inst : DFFRPQ1 port map( D => n164, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_2_port);
   arx_r2_reg_reg_2_inst : DFFRPQ1 port map( D => n144, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_2_port);
   arx_r3_reg_reg_2_inst : DFFRPQ1 port map( D => n159, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_2_port);
   arx_d2_reg_reg_12_inst : DFERPQ1 port map( D => arx_d1_reg_12_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => 
                           arx_d2_reg_12_port);
   arx_d2_reg_reg_13_inst : DFERPQ1 port map( D => arx_d1_reg_13_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => 
                           arx_d2_reg_13_port);
   arx_r1_reg_reg_0_inst : DFFRPQ1 port map( D => n162, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_0_port);
   arx_r2_reg_reg_0_inst : DFFRPQ1 port map( D => n146, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_0_port);
   arx_r1_reg_reg_1_inst : DFFRPQ1 port map( D => n163, CK => clock, RB => 
                           resetn, Q => arx_r1_reg_1_port);
   arx_r3_reg_reg_0_inst : DFFRPQ1 port map( D => n161, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_0_port);
   arx_r4_reg_reg_1_inst : DFERPQ1 port map( D => m3_out_1_port, CEB => n1100, 
                           CK => clock, RB => resetn, Q => arx_r4_reg_1_port);
   arx_d2_reg_reg_11_inst : DFERPQ1 port map( D => arx_d1_reg_11_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => 
                           arx_d2_reg_11_port);
   arx_r2_reg_reg_1_inst : DFFRPQ1 port map( D => n145, CK => clock, RB => 
                           resetn, Q => arx_r2_reg_1_port);
   arx_r3_reg_reg_1_inst : DFFRPQ1 port map( D => n160, CK => clock, RB => 
                           resetn, Q => arx_r3_reg_1_port);
   arx_d2_reg_reg_10_inst : DFERPQ1 port map( D => arx_d1_reg_10_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => 
                           arx_d2_reg_10_port);
   arx_d2_reg_reg_7_inst : DFERPQ1 port map( D => arx_d1_reg_7_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => 
                           arx_d2_reg_7_port);
   arx_d2_reg_reg_8_inst : DFERPQ1 port map( D => arx_d1_reg_8_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => 
                           arx_d2_reg_8_port);
   arx_d2_reg_reg_9_inst : DFERPQ1 port map( D => arx_d1_reg_9_port, CEB => 
                           n178, CK => clock, RB => resetn, Q => 
                           arx_d2_reg_9_port);
   arx_state_reg_reg_1_inst : DFFRPQ1 port map( D => n193, CK => clock, RB => 
                           resetn, Q => arx_state_reg_1_port);
   arx_state_reg_reg_0_inst : DFFRPQ1 port map( D => state_0_port, CK => clock,
                           RB => resetn, Q => arx_state_reg_0_port);
   arx_o1_reg_reg_7_inst : DFERPQ1 port map( D => a2_out_7_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => data_out(7));
   arx_o1_reg_reg_0_inst : DFERPQ1 port map( D => a2_out_0_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => data_out(0));
   arx_o1_reg_reg_1_inst : DFERPQ1 port map( D => a2_out_1_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => data_out(1));
   arx_o1_reg_reg_2_inst : DFERPQ1 port map( D => a2_out_2_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => data_out(2));
   arx_o1_reg_reg_3_inst : DFERPQ1 port map( D => a2_out_3_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => data_out(3));
   arx_o1_reg_reg_4_inst : DFERPQ1 port map( D => a2_out_4_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => data_out(4));
   arx_o1_reg_reg_5_inst : DFERPQ1 port map( D => a2_out_5_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => data_out(5));
   arx_o1_reg_reg_6_inst : DFERPQ1 port map( D => a2_out_6_port, CEB => n178, 
                           CK => clock, RB => resetn, Q => data_out(6));
   U249 : INVBD2 port map( A => arx_d2_reg_14_port, Z => n187);
   U250 : INVBD2 port map( A => arx_d2_reg_13_port, Z => n185);
   U251 : INVBD2 port map( A => arx_d2_reg_12_port, Z => n186);
   U252 : INVBD2 port map( A => arx_d2_reg_11_port, Z => n184);
   U253 : INVBD2 port map( A => arx_d2_reg_10_port, Z => n182);
   U254 : INVBD2 port map( A => arx_d2_reg_9_port, Z => n180);
   U255 : INVBD2 port map( A => arx_d2_reg_8_port, Z => n181);
   U256 : INVBD2 port map( A => arx_d2_reg_7_port, Z => n183);
   U257 : NOR2D2 port map( A1 => n231, A2 => n179, Z => a2_in_r_0_port);
   U258 : NOR2D2 port map( A1 => n202, A2 => arx_state_reg_1_port, Z => n177);
   U259 : OR2D1 port map( A1 => n177, A2 => state_0_port, Z => n178);
   U260 : NAN2D1 port map( A1 => arx_state_reg_0_port, A2 => 
                           arx_state_reg_1_port, Z => n179);
   U261 : INVD1 port map( A => n191, Z => n193);
   U262 : INVD1 port map( A => n192, Z => n191);
   U263 : INVD1 port map( A => n101, Z => n192);
   U264 : NAN2D1 port map( A1 => n193, A2 => n188, Z => n1100);
   U265 : INVD1 port map( A => m5_in_l_0, Z => n194);
   U266 : NOR2M1D1 port map( A1 => n179, A2 => n190, Z => n130);
   U267 : INVD1 port map( A => n189, Z => n188);
   U268 : NOR2D1 port map( A1 => n177, A2 => n190, Z => n101);
   U269 : NAN2D1 port map( A1 => n101, A2 => n179, Z => n127);
   U270 : NAN2M1D1 port map( A1 => n177, A2 => n129, Z => m5_in_l_0);
   U271 : NOR2D1 port map( A1 => n130, A2 => n216, Z => a2_in_l_1_port);
   U272 : NOR2D1 port map( A1 => n130, A2 => n217, Z => a2_in_l_0_port);
   U273 : INVD1 port map( A => n1110, Z => n190);
   U274 : NOR2D1 port map( A1 => n188, A2 => n224, Z => a1_in_l_0_port);
   U275 : NOR2D1 port map( A1 => n188, A2 => n218, Z => a1_in_l_6_port);
   U276 : NOR2D1 port map( A1 => n188, A2 => n222, Z => a1_in_l_2_port);
   U277 : NOR2D1 port map( A1 => n188, A2 => n221, Z => a1_in_l_3_port);
   U278 : NOR2D1 port map( A1 => n188, A2 => n220, Z => a1_in_l_4_port);
   U279 : INVD1 port map( A => n1110, Z => n189);
   U280 : NOR2D1 port map( A1 => n194, A2 => n248, Z => m2_in_r_0_port);
   U281 : NOR2D1 port map( A1 => n194, A2 => n201, Z => m2_in_r_1_port);
   U282 : NOR2D1 port map( A1 => n188, A2 => n223, Z => a1_in_l_1_port);
   U283 : NOR2D1 port map( A1 => n194, A2 => n200, Z => m2_in_r_2_port);
   U284 : NOR2D1 port map( A1 => n194, A2 => n199, Z => m2_in_r_3_port);
   U285 : NOR2D1 port map( A1 => n191, A2 => n198, Z => m1_in_r_4_port);
   U286 : NOR2D1 port map( A1 => n191, A2 => n199, Z => m1_in_r_3_port);
   U287 : NOR2D1 port map( A1 => n191, A2 => n248, Z => m1_in_r_0_port);
   U288 : NOR2D1 port map( A1 => n191, A2 => n201, Z => m1_in_r_1_port);
   U289 : NOR2D1 port map( A1 => n191, A2 => n200, Z => m1_in_r_2_port);
   U290 : NOR2D1 port map( A1 => n191, A2 => n197, Z => m1_in_r_5_port);
   U291 : NOR2D1 port map( A1 => n130, A2 => n212, Z => a2_in_l_5_port);
   U292 : NOR2D1 port map( A1 => n194, A2 => n198, Z => m2_in_r_4_port);
   U293 : NOR2D1 port map( A1 => n194, A2 => n196, Z => m2_in_r_6_port);
   U294 : NOR2D1 port map( A1 => n194, A2 => n197, Z => m2_in_r_5_port);
   U295 : NOR2D1 port map( A1 => n101, A2 => n196, Z => m1_in_r_6_port);
   U296 : NOR2D1 port map( A1 => n101, A2 => n195, Z => m1_in_r_7_port);
   U297 : NOR2D1 port map( A1 => n188, A2 => n219, Z => a1_in_l_5_port);
   U298 : NOR2D1 port map( A1 => n194, A2 => n195, Z => m2_in_r_7_port);
   U299 : NOR2D1 port map( A1 => n130, A2 => n203, Z => a2_in_l_14_port);
   U300 : NAN2D1 port map( A1 => n188, A2 => n129, Z => state_0_port);
   U301 : INVD1 port map( A => arx_state_reg_0_port, Z => n202);
   U302 : NOR2D1 port map( A1 => n180, A2 => n194, Z => m4_in_r_2_port);
   U303 : NOR2D1 port map( A1 => n181, A2 => n194, Z => m4_in_r_1_port);
   U304 : NOR2D1 port map( A1 => n182, A2 => n194, Z => m4_in_r_3_port);
   U305 : NOR2D1 port map( A1 => n183, A2 => n194, Z => m4_in_r_0_port);
   U306 : NAN2M1D1 port map( A1 => arx_state_reg_1_port, A2 => n202, Z => n129)
                           ;
   U307 : NOR2D1 port map( A1 => n130, A2 => n211, Z => a2_in_l_6_port);
   U308 : NOR2D1 port map( A1 => n130, A2 => n210, Z => a2_in_l_7_port);
   U309 : NOR2D1 port map( A1 => n130, A2 => n209, Z => a2_in_l_8_port);
   U310 : NOR2D1 port map( A1 => n130, A2 => n208, Z => a2_in_l_9_port);
   U311 : NOR2D1 port map( A1 => n130, A2 => n207, Z => a2_in_l_10_port);
   U312 : NOR2D1 port map( A1 => n130, A2 => n206, Z => a2_in_l_11_port);
   U313 : NOR2D1 port map( A1 => n130, A2 => n205, Z => a2_in_l_12_port);
   U314 : NOR2D1 port map( A1 => n130, A2 => n204, Z => a2_in_l_13_port);
   U315 : NOR2D1 port map( A1 => n130, A2 => n215, Z => a2_in_l_2_port);
   U316 : NOR2D1 port map( A1 => n130, A2 => n214, Z => a2_in_l_3_port);
   U317 : NOR2D1 port map( A1 => n130, A2 => n213, Z => a2_in_l_4_port);
   U318 : NOR2D1 port map( A1 => n184, A2 => n194, Z => m4_in_r_4_port);
   U319 : NAN2D1 port map( A1 => arx_state_reg_1_port, A2 => n202, Z => n1110);
   U320 : NOR2D1 port map( A1 => n185, A2 => n194, Z => m4_in_r_6_port);
   U321 : NOR2D1 port map( A1 => n186, A2 => n194, Z => m4_in_r_5_port);
   U322 : AND2D1 port map( A1 => N48, A2 => m5_in_l_0, Z => m5_in_r_4_port);
   U323 : AND2D1 port map( A1 => N45, A2 => m5_in_l_0, Z => m5_in_r_1_port);
   U324 : AND2D1 port map( A1 => N46, A2 => m5_in_l_0, Z => m5_in_r_2_port);
   U325 : AND2D1 port map( A1 => N47, A2 => m5_in_l_0, Z => m5_in_r_3_port);
   U326 : AND2D1 port map( A1 => N44, A2 => m5_in_l_0, Z => m5_in_r_0_port);
   U327 : NOR2D1 port map( A1 => n187, A2 => n194, Z => m4_in_r_7_port);
   U328 : AND2D1 port map( A1 => N49, A2 => m5_in_l_0, Z => m5_in_r_5_port);
   U329 : AND2D1 port map( A1 => N50, A2 => m5_in_l_0, Z => m5_in_r_6_port);
   U330 : AND2D1 port map( A1 => N51, A2 => m5_in_l_0, Z => m5_in_r_7_port);
   U331 : INVD1 port map( A => arx_r3_reg_1_port, Z => n230);
   U332 : INVD1 port map( A => arx_r2_reg_1_port, Z => n223);
   U333 : INVD1 port map( A => arx_r3_reg_0_port, Z => n231);
   U334 : INVD1 port map( A => arx_r1_reg_1_port, Z => n216);
   U335 : INVD1 port map( A => arx_r2_reg_0_port, Z => n224);
   U336 : INVD1 port map( A => arx_r1_reg_0_port, Z => n217);
   U337 : INVD1 port map( A => arx_r3_reg_2_port, Z => n229);
   U338 : INVD1 port map( A => arx_r2_reg_2_port, Z => n222);
   U339 : INVD1 port map( A => arx_r1_reg_2_port, Z => n215);
   U340 : INVD1 port map( A => arx_d1_reg_7_port, Z => n248);
   U341 : INVD1 port map( A => arx_d1_reg_8_port, Z => n201);
   U342 : INVD1 port map( A => arx_d1_reg_9_port, Z => n200);
   U343 : INVD1 port map( A => arx_r3_reg_3_port, Z => n228);
   U344 : AO22D1 port map( A1 => m4_out_6_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_6_port, Z => n155);
   U345 : INVD1 port map( A => arx_r2_reg_3_port, Z => n221);
   U346 : INVD1 port map( A => arx_r1_reg_3_port, Z => n214);
   U347 : AO22D1 port map( A1 => m2_out_6_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_6_port, Z => n140);
   U348 : INVD1 port map( A => arx_r3_reg_4_port, Z => n227);
   U349 : INVD1 port map( A => arx_r2_reg_4_port, Z => n220);
   U350 : INVD1 port map( A => arx_d1_reg_10_port, Z => n199);
   U351 : INVD1 port map( A => arx_r1_reg_4_port, Z => n213);
   U352 : AO22D1 port map( A1 => m4_out_5_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_5_port, Z => n156);
   U353 : INVD1 port map( A => arx_d1_reg_11_port, Z => n198);
   U354 : INVD1 port map( A => arx_r3_reg_5_port, Z => n226);
   U355 : INVD1 port map( A => arx_r2_reg_5_port, Z => n219);
   U356 : AO22D1 port map( A1 => m2_out_5_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_5_port, Z => n141);
   U357 : INVD1 port map( A => arx_r1_reg_5_port, Z => n212);
   U358 : INVD1 port map( A => arx_r3_reg_6_port, Z => n225);
   U359 : AO22D1 port map( A1 => m4_out_4_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_4_port, Z => n157);
   U360 : INVD1 port map( A => arx_d1_reg_12_port, Z => n197);
   U361 : INVD1 port map( A => arx_r2_reg_6_port, Z => n218);
   U362 : INVD1 port map( A => arx_r1_reg_6_port, Z => n211);
   U363 : INVD1 port map( A => arx_d1_reg_13_port, Z => n196);
   U364 : AO22D1 port map( A1 => m2_out_4_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_4_port, Z => n142);
   U365 : INVD1 port map( A => arx_d1_reg_14_port, Z => n195);
   U366 : AO22D1 port map( A1 => m4_out_3_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_3_port, Z => n158);
   U367 : INVD1 port map( A => arx_r3_reg_7_port, Z => n232);
   U368 : INVD1 port map( A => arx_r2_reg_7_port, Z => n240);
   U369 : INVD1 port map( A => arx_r1_reg_7_port, Z => n210);
   U370 : AO22D1 port map( A1 => m2_out_3_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_3_port, Z => n143);
   U371 : INVD1 port map( A => arx_r3_reg_8_port, Z => n233);
   U372 : INVD1 port map( A => arx_r2_reg_8_port, Z => n241);
   U373 : AO22D1 port map( A1 => m4_out_2_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_2_port, Z => n159);
   U374 : INVD1 port map( A => arx_r1_reg_8_port, Z => n209);
   U375 : AO22D1 port map( A1 => m2_out_2_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_2_port, Z => n144);
   U376 : INVD1 port map( A => arx_r3_reg_9_port, Z => n234);
   U377 : INVD1 port map( A => arx_r2_reg_9_port, Z => n242);
   U378 : INVD1 port map( A => arx_r1_reg_9_port, Z => n208);
   U379 : AO22D1 port map( A1 => m4_out_1_port, A2 => n177, B1 => n101, B2 => 
                           arx_r3_reg_1_port, Z => n160);
   U380 : AO22D1 port map( A1 => m2_out_1_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_1_port, Z => n145);
   U381 : INVD1 port map( A => arx_r3_reg_10_port, Z => n235);
   U382 : INVD1 port map( A => arx_r2_reg_10_port, Z => n243);
   U383 : INVD1 port map( A => arx_r1_reg_10_port, Z => n207);
   U384 : AO22D1 port map( A1 => m2_out_0_port, A2 => n177, B1 => n101, B2 => 
                           arx_r2_reg_0_port, Z => n146);
   U385 : AO22D1 port map( A1 => m4_out_0_port, A2 => n177, B1 => n191, B2 => 
                           arx_r3_reg_0_port, Z => n161);
   U386 : INVD1 port map( A => arx_r3_reg_11_port, Z => n236);
   U387 : INVD1 port map( A => arx_r2_reg_11_port, Z => n244);
   U388 : INVD1 port map( A => arx_r1_reg_11_port, Z => n206);
   U389 : INVD1 port map( A => arx_r3_reg_12_port, Z => n237);
   U390 : INVD1 port map( A => arx_r2_reg_12_port, Z => n245);
   U391 : INVD1 port map( A => arx_r1_reg_12_port, Z => n205);
   U392 : INVD1 port map( A => arx_r3_reg_13_port, Z => n238);
   U393 : INVD1 port map( A => arx_r2_reg_13_port, Z => n246);
   U394 : INVD1 port map( A => arx_r1_reg_13_port, Z => n204);
   U395 : INVD1 port map( A => arx_r3_reg_14_port, Z => n239);
   U396 : INVD1 port map( A => arx_r2_reg_14_port, Z => n247);
   U397 : INVD1 port map( A => arx_r1_reg_14_port, Z => n203);
   U398 : TIELO port map( Z => net1801);
   U399 : EXOR2D1 port map( A1 => N114, A2 => add_416_C243_rn_carry_7_port, Z 
                           => a1_out_7_port);
   U400 : AND2D1 port map( A1 => add_416_C243_rn_carry_6_port, A2 => N113, Z =>
                           add_416_C243_rn_carry_7_port);
   U401 : EXOR2D1 port map( A1 => N113, A2 => add_416_C243_rn_carry_6_port, Z 
                           => a1_out_6_port);
   U402 : AND2D1 port map( A1 => add_416_C243_rn_carry_5_port, A2 => N112, Z =>
                           add_416_C243_rn_carry_6_port);
   U403 : EXOR2D1 port map( A1 => N112, A2 => add_416_C243_rn_carry_5_port, Z 
                           => a1_out_5_port);
   U404 : AND2D1 port map( A1 => add_416_C243_rn_carry_4_port, A2 => N111, Z =>
                           add_416_C243_rn_carry_5_port);
   U405 : EXOR2D1 port map( A1 => N111, A2 => add_416_C243_rn_carry_4_port, Z 
                           => a1_out_4_port);
   U406 : AND2D1 port map( A1 => add_416_C243_rn_carry_3_port, A2 => N110, Z =>
                           add_416_C243_rn_carry_4_port);
   U407 : EXOR2D1 port map( A1 => N110, A2 => add_416_C243_rn_carry_3_port, Z 
                           => a1_out_3_port);
   U408 : AND2D1 port map( A1 => add_416_C243_rn_carry_2_port, A2 => N109, Z =>
                           add_416_C243_rn_carry_3_port);
   U409 : EXOR2D1 port map( A1 => N109, A2 => add_416_C243_rn_carry_2_port, Z 
                           => a1_out_2_port);
   U410 : AND2D1 port map( A1 => add_416_C243_rn_carry_1_port, A2 => N108, Z =>
                           add_416_C243_rn_carry_2_port);
   U411 : EXOR2D1 port map( A1 => N108, A2 => add_416_C243_rn_carry_1_port, Z 
                           => a1_out_1_port);
   U412 : AND2D1 port map( A1 => N107, A2 => N106, Z => 
                           add_416_C243_rn_carry_1_port);
   U413 : EXOR2D1 port map( A1 => N106, A2 => N107, Z => a1_out_0_port);
   U414 : EXOR2D1 port map( A1 => N123, A2 => add_416_C244_rn_carry_7_port, Z 
                           => a2_out_7_port);
   U415 : AND2D1 port map( A1 => add_416_C244_rn_carry_6_port, A2 => N122, Z =>
                           add_416_C244_rn_carry_7_port);
   U416 : EXOR2D1 port map( A1 => N122, A2 => add_416_C244_rn_carry_6_port, Z 
                           => a2_out_6_port);
   U417 : AND2D1 port map( A1 => add_416_C244_rn_carry_5_port, A2 => N121, Z =>
                           add_416_C244_rn_carry_6_port);
   U418 : EXOR2D1 port map( A1 => N121, A2 => add_416_C244_rn_carry_5_port, Z 
                           => a2_out_5_port);
   U419 : AND2D1 port map( A1 => add_416_C244_rn_carry_4_port, A2 => N120, Z =>
                           add_416_C244_rn_carry_5_port);
   U420 : EXOR2D1 port map( A1 => N120, A2 => add_416_C244_rn_carry_4_port, Z 
                           => a2_out_4_port);
   U421 : AND2D1 port map( A1 => add_416_C244_rn_carry_3_port, A2 => N119, Z =>
                           add_416_C244_rn_carry_4_port);
   U422 : EXOR2D1 port map( A1 => N119, A2 => add_416_C244_rn_carry_3_port, Z 
                           => a2_out_3_port);
   U423 : AND2D1 port map( A1 => add_416_C244_rn_carry_2_port, A2 => N118, Z =>
                           add_416_C244_rn_carry_3_port);
   U424 : EXOR2D1 port map( A1 => N118, A2 => add_416_C244_rn_carry_2_port, Z 
                           => a2_out_2_port);
   U425 : AND2D1 port map( A1 => add_416_C244_rn_carry_1_port, A2 => N117, Z =>
                           add_416_C244_rn_carry_2_port);
   U426 : EXOR2D1 port map( A1 => N117, A2 => add_416_C244_rn_carry_1_port, Z 
                           => a2_out_1_port);
   U427 : AND2D1 port map( A1 => N116, A2 => N115, Z => 
                           add_416_C244_rn_carry_1_port);
   U428 : EXOR2D1 port map( A1 => N115, A2 => N116, Z => a2_out_0_port);

end hier_rtl_none_10;
