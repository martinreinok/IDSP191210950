--
-- MAP7_overlapped_std
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.arx_numeric.all;

entity MAP7_overlapped_std is
   port(
      clock : in std_logic;
      resetn : in std_logic;
      data_in : in std_logic_vector(7 downto 0);
      data1_out : out std_logic_vector(7 downto 0)
   );
end MAP7_overlapped_std;

architecture rtl of MAP7_overlapped_std is
   component MAP7_overlapped
      port (
         clock : in std_logic;
         resetn : in std_logic;
         data_in : in signed(7 downto 0);
         data1_out : out signed(7 downto 0)
      );
   end component;

   signal arx_data_in : signed(7 downto 0);
   signal arx_data1_out : signed(7 downto 0);
begin

   MAP7_overlapped_inst : MAP7_overlapped
      port map (
         clock => clock,
         resetn => resetn,
         data_in => arx_data_in,
         data1_out => arx_data1_out
      );

   arx_data_in <= signed(data_in);
   data1_out <= std_logic_vector(arx_data1_out);
end rtl;

--
-- MAP7_overlapped
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.arx_numeric.all;

entity MAP7_overlapped is
   port(
      clock : in std_logic;
      resetn : in std_logic;
      data_in : in signed(7 downto 0);
      data1_out : out signed(7 downto 0)
   );
end MAP7_overlapped;

architecture rtl of MAP7_overlapped is
   type T_state is (T_state_cycle0, T_state_cycle1, T_state_cycle2, T_state_cycle3);

   constant arx_i1_reset : signed(7 downto 0) := "00000000";
   constant arx_o1_reset : signed(7 downto 0) := "00000000";
   constant arx_r1_reset : signed(15 downto 0) := "0000000000000000";
   constant arx_r2_reset : signed(15 downto 0) := "0000000000000000";
   constant arx_r3_reset : signed(15 downto 0) := "0000000000000000";
   constant arx_r4_reset : signed(15 downto 0) := "0000000000000000";
   constant arx_d1_reset : signed(15 downto 0) := "0000000000000000";
   constant arx_d2_reset : signed(15 downto 0) := "0000000000000000";
   constant arx_state_reset : T_state := T_state_cycle0;

   signal arx_i1_reg, arx_i1_nxt : signed(7 downto 0);
   signal arx_o1_reg, arx_o1_nxt : signed(7 downto 0);
   signal arx_r1_reg, arx_r1_nxt : signed(15 downto 0);
   signal arx_r2_reg, arx_r2_nxt : signed(15 downto 0);
   signal arx_r3_reg, arx_r3_nxt : signed(15 downto 0);
   signal arx_r4_reg, arx_r4_nxt : signed(15 downto 0);
   signal arx_d1_reg, arx_d1_nxt : signed(15 downto 0);
   signal arx_d2_reg, arx_d2_nxt : signed(15 downto 0);
   signal arx_state_reg, arx_state_nxt : T_state;
begin

   registers : process (resetn, clock)
   begin
      if resetn = '0' then
         arx_i1_reg <= arx_i1_reset;
         arx_o1_reg <= arx_o1_reset;
         arx_r1_reg <= arx_r1_reset;
         arx_r2_reg <= arx_r2_reset;
         arx_r3_reg <= arx_r3_reset;
         arx_r4_reg <= arx_r4_reset;
         arx_d1_reg <= arx_d1_reset;
         arx_d2_reg <= arx_d2_reset;
         arx_state_reg <= arx_state_reset;
      elsif rising_edge(clock) then
         arx_i1_reg <= arx_i1_nxt;
         arx_o1_reg <= arx_o1_nxt;
         arx_r1_reg <= arx_r1_nxt;
         arx_r2_reg <= arx_r2_nxt;
         arx_r3_reg <= arx_r3_nxt;
         arx_r4_reg <= arx_r4_nxt;
         arx_d1_reg <= arx_d1_nxt;
         arx_d2_reg <= arx_d2_nxt;
         arx_state_reg <= arx_state_nxt;
      end if;
   end process registers;

   update : process (data_in, arx_i1_reg, arx_o1_reg, arx_r1_reg, arx_r2_reg, arx_r3_reg, arx_r4_reg, arx_d1_reg, arx_d2_reg, arx_state_reg)
      variable m1_in_l : signed(7 downto 0); -- reads=1, writes=4
      variable m1_in_r : signed(7 downto 0); -- reads=1, writes=4
      variable m1_out : signed(15 downto 0); -- reads=2, writes=1
      variable m2_in_l : signed(7 downto 0); -- reads=1, writes=4
      variable m2_in_r : signed(7 downto 0); -- reads=1, writes=4
      variable m2_out : signed(15 downto 0); -- reads=2, writes=1
      variable m3_in_l : signed(7 downto 0); -- reads=1, writes=2
      variable m3_in_r : signed(7 downto 0); -- reads=1, writes=2
      variable m3_out : signed(15 downto 0); -- reads=1, writes=1
      variable a1_in_l : signed(15 downto 0); -- reads=1, writes=3
      variable a1_in_r : signed(15 downto 0); -- reads=1, writes=3
      variable a1_out : signed(7 downto 0); -- reads=3, writes=1
      variable a2_in_l : signed(15 downto 0); -- reads=1, writes=1
      variable a2_in_r : signed(15 downto 0); -- reads=1, writes=1
      variable a2_out : signed(7 downto 0); -- reads=1, writes=1
      variable b2 : signed(7 downto 0); -- reads=2, writes=1
      variable b1 : signed(7 downto 0); -- reads=2, writes=1
      variable b0 : signed(7 downto 0); -- reads=2, writes=1
      variable a2 : signed(7 downto 0); -- reads=2, writes=1
      variable a1 : signed(7 downto 0); -- reads=2, writes=1
      variable i1 : signed(7 downto 0); -- reads=1, writes=1
      variable o1 : signed(7 downto 0); -- reads=1, writes=1
      variable r1 : signed(15 downto 0); -- reads=2, writes=2
      variable r2 : signed(15 downto 0); -- reads=3, writes=3
      variable r3 : signed(15 downto 0); -- reads=1, writes=1
      variable r4 : signed(15 downto 0); -- reads=1, writes=1
      variable d1 : signed(15 downto 0); -- reads=7, writes=1
      variable d2 : signed(15 downto 0); -- reads=4, writes=1
      variable state : T_state; -- reads=3, writes=4
   begin
      --initialize variables and outports
      m1_in_l := to_signed(0, 8);
      m1_in_r := to_signed(0, 8);
      m1_out := to_signed(0, 16);
      m2_in_l := to_signed(0, 8);
      m2_in_r := to_signed(0, 8);
      m2_out := to_signed(0, 16);
      m3_in_l := to_signed(0, 8);
      m3_in_r := to_signed(0, 8);
      m3_out := to_signed(0, 16);
      a1_in_l := to_signed(0, 16);
      a1_in_r := to_signed(0, 16);
      a1_out := to_signed(0, 8);
      a2_in_l := to_signed(0, 16);
      a2_in_r := to_signed(0, 16);
      a2_out := to_signed(0, 8);
      b2 := to_signed(0, 8);
      b1 := to_signed(0, 8);
      b0 := to_signed(0, 8);
      a2 := to_signed(0, 8);
      a1 := to_signed(0, 8);
      data1_out <= to_signed(0, 8);
      --copy register values to local variables
      i1 := arx_i1_reg;
      o1 := arx_o1_reg;
      r1 := arx_r1_reg;
      r2 := arx_r2_reg;
      r3 := arx_r3_reg;
      r4 := arx_r4_reg;
      d1 := arx_d1_reg;
      d2 := arx_d2_reg;
      state := arx_state_reg;
      --read from component outports
      --update outputs and register values
      b2 := "00111001";
      b1 := "10011010";
      b0 := "00111001";
      a2 := "11001111";
      a1 := "01000011";
      case arx_state_reg is
         when T_state_cycle0 =>
            m1_in_l := b1;
            m1_in_r := arx_wrap(arx_round(arx_d1_reg, 7), 1);
            m2_in_l := b2;
            m2_in_r := arx_wrap(arx_round(arx_d2_reg, 7), 1);
         when T_state_cycle1 =>
            m1_in_l := b1;
            m1_in_r := arx_wrap(arx_round(arx_d1_reg, 7), 1);
            m2_in_l := b2;
            m2_in_r := arx_wrap(arx_round(arx_d2_reg, 7), 1);
         when T_state_cycle2 =>
            m1_in_l := a1;
            m1_in_r := arx_wrap(arx_round(arx_d1_reg, 7), 1);
            m2_in_l := a2;
            m2_in_r := arx_wrap(arx_round(arx_d2_reg, 7), 1);
            m3_in_l := b0;
            m3_in_r := arx_wrap(arx_round(arx_d1_reg, 7), 1);
         when T_state_cycle3 =>
            m1_in_l := a1;
            m1_in_r := arx_wrap(arx_round(arx_d1_reg, 7), 1);
            m2_in_l := a2;
            m2_in_r := arx_wrap(arx_round(arx_d2_reg, 7), 1);
            m3_in_l := b0;
            m3_in_r := arx_wrap(arx_round(arx_d1_reg, 7), 1);
      end case;
      case arx_state_reg is
         when T_state_cycle0 =>
            a1_in_l := arx_r1_reg;
            a1_in_r := arx_r2_reg;
            a2_in_l := arx_r3_reg;
            a2_in_r := arx_r4_reg;
         when T_state_cycle1 =>
            a1_in_l := arx_msb_extend(arx_lsb_extend(arx_i1_reg, 7), 1);
            a1_in_r := arx_r2_reg;
         when T_state_cycle2 =>
            a1_in_l := arx_r1_reg;
            a1_in_r := arx_r2_reg;
         when T_state_cycle3 =>
      end case;
      m1_out := (m1_in_l * m1_in_r);
      m2_out := (m2_in_l * m2_in_r);
      m3_out := (m3_in_l * m3_in_r);
      a1_out := arx_wrap(arx_round((arx_msb_extend(a1_in_l, 1) + arx_msb_extend(a1_in_r, 1)), 7), 2);
      a2_out := arx_wrap(arx_round((arx_msb_extend(a2_in_l, 1) + arx_msb_extend(a2_in_r, 1)), 7), 2);
      case arx_state_reg is
         when T_state_cycle0 =>
            state := T_state_cycle1;
            i1 := data_in;
            r2 := arx_msb_extend(arx_lsb_extend(a1_out, 7), 1);
            o1 := a2_out;
         when T_state_cycle1 =>
            state := T_state_cycle2;
            r1 := m1_out;
            r2 := m2_out;
            d2 := arx_d1_reg;
            d1 := arx_msb_extend(arx_lsb_extend(a1_out, 7), 1);
         when T_state_cycle2 =>
            state := T_state_cycle3;
            r3 := arx_msb_extend(arx_lsb_extend(a1_out, 7), 1);
         when T_state_cycle3 =>
            state := T_state_cycle0;
            r1 := m1_out;
            r2 := m2_out;
            r4 := m3_out;
      end case;
      data1_out <= arx_o1_reg;
      --write to component inports
      --copy local variables to next register values
      arx_i1_nxt <= i1;
      arx_o1_nxt <= o1;
      arx_r1_nxt <= r1;
      arx_r2_nxt <= r2;
      arx_r3_nxt <= r3;
      arx_r4_nxt <= r4;
      arx_d1_nxt <= d1;
      arx_d2_nxt <= d2;
      arx_state_nxt <= state;
   end process update;
end rtl;

