
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_gfsk is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_gfsk;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_gfsk.all;

architecture flat_structure_none_10 of gfsk is

   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI31M10D1
      port( A1, A2, A3, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   component NOR4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI31D1
      port( A1, A2, A3, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22M20D1
      port( B1, B2, A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN4D1
      port( A1, A2, A3, A4 : in std_logic;  Z : out std_logic);
   end component;
   
   component BUFD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component EXNOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component TIEHI
      port( Z : out std_logic);
   end component;
   
   signal n_Logic1, n_Logic0, slicer_out_port, clk4, mixer_out_i_11_port, 
      mixer_out_i_10_port, mixer_out_i_9_port, mixer_out_i_8_port, 
      mixer_out_i_7_port, mixer_out_i_6_port, mixer_out_i_5_port, 
      mixer_out_i_4_port, mixer_out_i_3_port, mixer_out_i_2_port, 
      mixer_out_i_1_port, mixer_out_i_0_port, mixer_out_q_11_port, 
      mixer_out_q_10_port, mixer_out_q_9_port, mixer_out_q_8_port, 
      mixer_out_q_7_port, mixer_out_q_6_port, mixer_out_q_5_port, 
      mixer_out_q_4_port, mixer_out_q_3_port, mixer_out_q_2_port, 
      mixer_out_q_1_port, mixer_out_q_0_port, filter_out_i_4_port, 
      filter_out_i_3_port, filter_out_i_2_port, filter_out_i_1_port, 
      filter_out_i_0_port, filter_out_q_4_port, filter_out_q_3_port, 
      filter_out_q_2_port, filter_out_q_1_port, filter_out_q_0_port, 
      demodulator_out_6_port, demodulator_out_5_port, demodulator_out_4_port, 
      demodulator_out_3_port, demodulator_out_2_port, demodulator_out_1_port, 
      demodulator_out_0_port, cg_n10, cg_N2, cg_N1, cg_counter_0_port, 
      cg_counter_1_port, mx_mixer_inst_n_1441, mx_mixer_inst_n_1440, 
      mx_mixer_inst_n_1439, mx_mixer_inst_n_1438, mx_mixer_inst_n_1437, 
      mx_mixer_inst_n_1436, mx_mixer_inst_n_1435, mx_mixer_inst_n_1434, 
      mx_mixer_inst_n_1433, mx_mixer_inst_n_1432, mx_mixer_inst_n_1431, 
      mx_mixer_inst_n_1430, mx_mixer_inst_n_1429, mx_mixer_inst_n_1428, 
      mx_mixer_inst_n88, mx_mixer_inst_n87, mx_mixer_inst_n86, 
      mx_mixer_inst_n85, mx_mixer_inst_n84, mx_mixer_inst_n83, 
      mx_mixer_inst_n82, mx_mixer_inst_n81, mx_mixer_inst_n80, 
      mx_mixer_inst_n79, mx_mixer_inst_n78, mx_mixer_inst_n77, 
      mx_mixer_inst_n76, mx_mixer_inst_n75, mx_mixer_inst_n74, 
      mx_mixer_inst_n73, mx_mixer_inst_n72, mx_mixer_inst_n71, 
      mx_mixer_inst_n70, mx_mixer_inst_n69, mx_mixer_inst_n680, 
      mx_mixer_inst_n670, mx_mixer_inst_n660, mx_mixer_inst_n650, 
      mx_mixer_inst_n640, mx_mixer_inst_n630, mx_mixer_inst_n620, 
      mx_mixer_inst_n610, mx_mixer_inst_n600, mx_mixer_inst_n590, 
      mx_mixer_inst_n580, mx_mixer_inst_n570, mx_mixer_inst_n560, 
      mx_mixer_inst_n550, mx_mixer_inst_n540, mx_mixer_inst_n530, 
      mx_mixer_inst_n520, mx_mixer_inst_n510, mx_mixer_inst_n500, 
      mx_mixer_inst_n490, mx_mixer_inst_n480, mx_mixer_inst_n470, 
      mx_mixer_inst_n460, mx_mixer_inst_n450, mx_mixer_inst_n440, 
      mx_mixer_inst_n430, mx_mixer_inst_n420, mx_mixer_inst_n410, 
      mx_mixer_inst_n400, mx_mixer_inst_n390, mx_mixer_inst_n380, 
      mx_mixer_inst_n370, mx_mixer_inst_n360, mx_mixer_inst_n350, 
      mx_mixer_inst_n340, mx_mixer_inst_n330, mx_mixer_inst_n32, 
      mx_mixer_inst_n31, mx_mixer_inst_n30, mx_mixer_inst_n29, 
      mx_mixer_inst_n28, mx_mixer_inst_n27, mx_mixer_inst_n26, 
      mx_mixer_inst_n25, mx_mixer_inst_n24, mx_mixer_inst_n23, 
      mx_mixer_inst_n22, mx_mixer_inst_n21, mx_mixer_inst_n20, 
      mx_mixer_inst_n19, mx_mixer_inst_n18, mx_mixer_inst_n17, 
      mx_mixer_inst_n16, mx_mixer_inst_n15, mx_mixer_inst_n14, 
      mx_mixer_inst_n13, mx_mixer_inst_n12, mx_mixer_inst_n11, 
      mx_mixer_inst_n10, mx_mixer_inst_n9, mx_mixer_inst_n8, mx_mixer_inst_n7, 
      mx_mixer_inst_n6, mx_mixer_inst_n5, mx_mixer_inst_n4, mx_mixer_inst_n3, 
      mx_mixer_inst_n2, mx_mixer_inst_n1, mx_mixer_inst_r377_carry_16_port, 
      mx_mixer_inst_r377_carry_15_port, mx_mixer_inst_r377_carry_14_port, 
      mx_mixer_inst_r377_carry_13_port, mx_mixer_inst_r377_carry_12_port, 
      mx_mixer_inst_r377_carry_11_port, mx_mixer_inst_r377_carry_10_port, 
      mx_mixer_inst_r377_carry_9_port, mx_mixer_inst_r377_carry_8_port, 
      mx_mixer_inst_N68, mx_mixer_inst_N67, mx_mixer_inst_N66, 
      mx_mixer_inst_N65, mx_mixer_inst_N64, mx_mixer_inst_N63, 
      mx_mixer_inst_N62, mx_mixer_inst_N61, mx_mixer_inst_N60, 
      mx_mixer_inst_N59, mx_mixer_inst_N58, mx_mixer_inst_N55, 
      mx_mixer_inst_N54, mx_mixer_inst_N53, mx_mixer_inst_N52, 
      mx_mixer_inst_N51, mx_mixer_inst_N50, mx_mixer_inst_N49, 
      mx_mixer_inst_N48, mx_mixer_inst_N47, mx_mixer_inst_N46, 
      mx_mixer_inst_N45, mx_mixer_inst_N44, mx_mixer_inst_N43, 
      mx_mixer_inst_N42, mx_mixer_inst_N41, mx_mixer_inst_N40, 
      mx_mixer_inst_N39, mx_mixer_inst_N38, mx_mixer_inst_N37, 
      mx_mixer_inst_N36, mx_mixer_inst_N35, mx_mixer_inst_N34, 
      mx_mixer_inst_N33, mx_mixer_inst_i_1_port, mx_mixer_inst_i_2_port, 
      mx_mixer_inst_arx_i_reg_0_port, mx_mixer_inst_arx_i_reg_1_port, 
      mx_mixer_inst_arx_i_reg_2_port, mx_mixer_inst_r375_n135, 
      mx_mixer_inst_r375_n134, mx_mixer_inst_r375_n133, mx_mixer_inst_r375_n132
      , mx_mixer_inst_r375_n131, mx_mixer_inst_r375_n130, 
      mx_mixer_inst_r375_n129, mx_mixer_inst_r375_n128, mx_mixer_inst_r375_n127
      , mx_mixer_inst_r375_n126, mx_mixer_inst_r375_n125, 
      mx_mixer_inst_r375_n124, mx_mixer_inst_r375_n123, mx_mixer_inst_r375_n122
      , mx_mixer_inst_r375_n121, mx_mixer_inst_r375_n120, 
      mx_mixer_inst_r375_n119, mx_mixer_inst_r375_n118, mx_mixer_inst_r375_n117
      , mx_mixer_inst_r375_n116, mx_mixer_inst_r375_n115, 
      mx_mixer_inst_r375_n114, mx_mixer_inst_r375_n113, mx_mixer_inst_r375_n53,
      mx_mixer_inst_r375_n52, mx_mixer_inst_r375_n51, mx_mixer_inst_r375_n50, 
      mx_mixer_inst_r375_n49, mx_mixer_inst_r375_n48, mx_mixer_inst_r375_n47, 
      mx_mixer_inst_r375_n46, mx_mixer_inst_r375_n45, mx_mixer_inst_r375_n44, 
      mx_mixer_inst_r375_n43, mx_mixer_inst_r375_n42, mx_mixer_inst_r375_n41, 
      mx_mixer_inst_r375_n40, mx_mixer_inst_r375_n39, mx_mixer_inst_r375_n38, 
      mx_mixer_inst_r375_n37, mx_mixer_inst_r375_n36, mx_mixer_inst_r375_n35, 
      mx_mixer_inst_r375_n34, mx_mixer_inst_r375_n33, mx_mixer_inst_r375_n32, 
      mx_mixer_inst_r375_n31, mx_mixer_inst_r375_n30, mx_mixer_inst_r375_n29, 
      mx_mixer_inst_r375_n28, mx_mixer_inst_r375_n27, mx_mixer_inst_r375_n26, 
      mx_mixer_inst_r375_n25, mx_mixer_inst_r375_n24, mx_mixer_inst_r375_n23, 
      mx_mixer_inst_r375_n22, mx_mixer_inst_r375_n21, mx_mixer_inst_r375_n20, 
      mx_mixer_inst_r375_n19, mx_mixer_inst_r375_n18, mx_mixer_inst_r375_n13, 
      mx_mixer_inst_r375_n12, mx_mixer_inst_r375_n11, mx_mixer_inst_r375_n10, 
      mx_mixer_inst_r375_n9, mx_mixer_inst_r375_n8, mx_mixer_inst_r375_n7, 
      mx_mixer_inst_r375_n6, mx_mixer_inst_r375_n5, mx_mixer_inst_r375_n4, 
      mx_mixer_inst_r375_n3, mx_mixer_inst_r375_n2, mx_mixer_inst_r376_n104, 
      mx_mixer_inst_r376_n103, mx_mixer_inst_r376_n102, mx_mixer_inst_r376_n101
      , mx_mixer_inst_r376_n100, mx_mixer_inst_r376_n99, mx_mixer_inst_r376_n98
      , mx_mixer_inst_r376_n97, mx_mixer_inst_r376_n96, mx_mixer_inst_r376_n95,
      mx_mixer_inst_r376_n94, mx_mixer_inst_r376_n52, mx_mixer_inst_r376_n51, 
      mx_mixer_inst_r376_n50, mx_mixer_inst_r376_n49, mx_mixer_inst_r376_n48, 
      mx_mixer_inst_r376_n47, mx_mixer_inst_r376_n46, mx_mixer_inst_r376_n45, 
      mx_mixer_inst_r376_n44, mx_mixer_inst_r376_n43, mx_mixer_inst_r376_n42, 
      mx_mixer_inst_r376_n41, mx_mixer_inst_r376_n40, mx_mixer_inst_r376_n39, 
      mx_mixer_inst_r376_n38, mx_mixer_inst_r376_n37, mx_mixer_inst_r376_n36, 
      mx_mixer_inst_r376_n35, mx_mixer_inst_r376_n34, mx_mixer_inst_r376_n33, 
      mx_mixer_inst_r376_n32, mx_mixer_inst_r376_n31, mx_mixer_inst_r376_n30, 
      mx_mixer_inst_r376_n29, mx_mixer_inst_r376_n28, mx_mixer_inst_r376_n27, 
      mx_mixer_inst_r376_n26, mx_mixer_inst_r376_n25, mx_mixer_inst_r376_n24, 
      mx_mixer_inst_r376_n23, mx_mixer_inst_r376_n22, mx_mixer_inst_r376_n21, 
      mx_mixer_inst_r376_n20, mx_mixer_inst_r376_n19, mx_mixer_inst_r376_n18, 
      mx_mixer_inst_r376_n17, mx_mixer_inst_r376_n16, mx_mixer_inst_r376_n15, 
      mx_mixer_inst_r376_n11, mx_mixer_inst_r376_n10, mx_mixer_inst_r376_n9, 
      mx_mixer_inst_r376_n8, mx_mixer_inst_r376_n7, mx_mixer_inst_r376_n6, 
      mx_mixer_inst_r376_n5, mx_mixer_inst_r376_n4, mx_mixer_inst_r376_n3, 
      mx_mixer_inst_r376_n2, lpf_filter_inst_lpf_i_n_1421, 
      lpf_filter_inst_lpf_i_n_1420, lpf_filter_inst_lpf_i_n_1419, 
      lpf_filter_inst_lpf_i_n_1418, lpf_filter_inst_lpf_i_n_1417, 
      lpf_filter_inst_lpf_i_n_1416, lpf_filter_inst_lpf_i_n_1415, 
      lpf_filter_inst_lpf_i_n_1414, lpf_filter_inst_lpf_i_n_1413, 
      lpf_filter_inst_lpf_i_n_1412, lpf_filter_inst_lpf_i_n_1411, 
      lpf_filter_inst_lpf_i_n_1410, lpf_filter_inst_lpf_i_n_1409, 
      lpf_filter_inst_lpf_i_n_1408, lpf_filter_inst_lpf_i_n_1407, 
      lpf_filter_inst_lpf_i_n_1406, lpf_filter_inst_lpf_i_n_1405, 
      lpf_filter_inst_lpf_i_n_1404, lpf_filter_inst_lpf_i_n_1403, 
      lpf_filter_inst_lpf_i_n_1402, lpf_filter_inst_lpf_i_n_1401, 
      lpf_filter_inst_lpf_i_n_1400, lpf_filter_inst_lpf_i_n_1399, 
      lpf_filter_inst_lpf_i_n_1398, lpf_filter_inst_lpf_i_n_1397, 
      lpf_filter_inst_lpf_i_n_1396, lpf_filter_inst_lpf_i_n_1395, 
      lpf_filter_inst_lpf_i_n_1394, lpf_filter_inst_lpf_i_n_1393, 
      lpf_filter_inst_lpf_i_n_1392, lpf_filter_inst_lpf_i_n_1391, 
      lpf_filter_inst_lpf_i_n_1390, lpf_filter_inst_lpf_i_n_1389, 
      lpf_filter_inst_lpf_i_n_1388, lpf_filter_inst_lpf_i_n_1387, 
      lpf_filter_inst_lpf_i_n_1386, lpf_filter_inst_lpf_i_n_1385, 
      lpf_filter_inst_lpf_i_n_1384, lpf_filter_inst_lpf_i_n_1383, 
      lpf_filter_inst_lpf_i_n_1382, lpf_filter_inst_lpf_i_n_1381, 
      lpf_filter_inst_lpf_i_n_1380, lpf_filter_inst_lpf_i_n_1379, 
      lpf_filter_inst_lpf_i_n_1378, lpf_filter_inst_lpf_i_n_1377, 
      lpf_filter_inst_lpf_i_n_1376, lpf_filter_inst_lpf_i_n_1375, 
      lpf_filter_inst_lpf_i_n_1374, lpf_filter_inst_lpf_i_n_1373, 
      lpf_filter_inst_lpf_i_n_1372, lpf_filter_inst_lpf_i_n194, 
      lpf_filter_inst_lpf_i_n193, lpf_filter_inst_lpf_i_n192, 
      lpf_filter_inst_lpf_i_n191, lpf_filter_inst_lpf_i_n190, 
      lpf_filter_inst_lpf_i_n189, lpf_filter_inst_lpf_i_n188, 
      lpf_filter_inst_lpf_i_n187, lpf_filter_inst_lpf_i_n186, 
      lpf_filter_inst_lpf_i_n185, lpf_filter_inst_lpf_i_n184, 
      lpf_filter_inst_lpf_i_n183, lpf_filter_inst_lpf_i_n182, 
      lpf_filter_inst_lpf_i_n181, lpf_filter_inst_lpf_i_n180, 
      lpf_filter_inst_lpf_i_n179, lpf_filter_inst_lpf_i_n178, 
      lpf_filter_inst_lpf_i_n177, lpf_filter_inst_lpf_i_n176, 
      lpf_filter_inst_lpf_i_n175, lpf_filter_inst_lpf_i_n174, 
      lpf_filter_inst_lpf_i_n173, lpf_filter_inst_lpf_i_n172, 
      lpf_filter_inst_lpf_i_n171, lpf_filter_inst_lpf_i_n170, 
      lpf_filter_inst_lpf_i_n169, lpf_filter_inst_lpf_i_n168, 
      lpf_filter_inst_lpf_i_n167, lpf_filter_inst_lpf_i_n166, 
      lpf_filter_inst_lpf_i_n165, lpf_filter_inst_lpf_i_n164, 
      lpf_filter_inst_lpf_i_n163, lpf_filter_inst_lpf_i_n162, 
      lpf_filter_inst_lpf_i_n161, lpf_filter_inst_lpf_i_n160, 
      lpf_filter_inst_lpf_i_n159, lpf_filter_inst_lpf_i_n157, 
      lpf_filter_inst_lpf_i_n156, lpf_filter_inst_lpf_i_n155, 
      lpf_filter_inst_lpf_i_n154, lpf_filter_inst_lpf_i_n153, 
      lpf_filter_inst_lpf_i_n152, lpf_filter_inst_lpf_i_n151, 
      lpf_filter_inst_lpf_i_n150, lpf_filter_inst_lpf_i_n149, 
      lpf_filter_inst_lpf_i_n148, lpf_filter_inst_lpf_i_n147, 
      lpf_filter_inst_lpf_i_n146, lpf_filter_inst_lpf_i_n145, 
      lpf_filter_inst_lpf_i_n144, lpf_filter_inst_lpf_i_n143, 
      lpf_filter_inst_lpf_i_n142, lpf_filter_inst_lpf_i_n141, 
      lpf_filter_inst_lpf_i_n140, lpf_filter_inst_lpf_i_n139, 
      lpf_filter_inst_lpf_i_n138, lpf_filter_inst_lpf_i_n137, 
      lpf_filter_inst_lpf_i_n136, lpf_filter_inst_lpf_i_n135, 
      lpf_filter_inst_lpf_i_n134, lpf_filter_inst_lpf_i_n133, 
      lpf_filter_inst_lpf_i_n132, lpf_filter_inst_lpf_i_n131, 
      lpf_filter_inst_lpf_i_n130, lpf_filter_inst_lpf_i_n129, 
      lpf_filter_inst_lpf_i_n128, lpf_filter_inst_lpf_i_n127, 
      lpf_filter_inst_lpf_i_n126, lpf_filter_inst_lpf_i_n125, 
      lpf_filter_inst_lpf_i_n124, lpf_filter_inst_lpf_i_n123, 
      lpf_filter_inst_lpf_i_n122, lpf_filter_inst_lpf_i_n121, 
      lpf_filter_inst_lpf_i_n120, lpf_filter_inst_lpf_i_n119, 
      lpf_filter_inst_lpf_i_n118, lpf_filter_inst_lpf_i_n117, 
      lpf_filter_inst_lpf_i_n116, lpf_filter_inst_lpf_i_n115, 
      lpf_filter_inst_lpf_i_n114, lpf_filter_inst_lpf_i_n113, 
      lpf_filter_inst_lpf_i_n112, lpf_filter_inst_lpf_i_n111, 
      lpf_filter_inst_lpf_i_n110, lpf_filter_inst_lpf_i_n109, 
      lpf_filter_inst_lpf_i_n108, lpf_filter_inst_lpf_i_n107, 
      lpf_filter_inst_lpf_i_n106, lpf_filter_inst_lpf_i_n105, 
      lpf_filter_inst_lpf_i_n104, lpf_filter_inst_lpf_i_n103, 
      lpf_filter_inst_lpf_i_n102, lpf_filter_inst_lpf_i_n101, 
      lpf_filter_inst_lpf_i_n100, lpf_filter_inst_lpf_i_n99, 
      lpf_filter_inst_lpf_i_n98, lpf_filter_inst_lpf_i_n97, 
      lpf_filter_inst_lpf_i_n96, lpf_filter_inst_lpf_i_n95, 
      lpf_filter_inst_lpf_i_n94, lpf_filter_inst_lpf_i_n92, 
      lpf_filter_inst_lpf_i_n91, lpf_filter_inst_lpf_i_n90, 
      lpf_filter_inst_lpf_i_n89, lpf_filter_inst_lpf_i_n88, 
      lpf_filter_inst_lpf_i_n87, lpf_filter_inst_lpf_i_n86, 
      lpf_filter_inst_lpf_i_n85, lpf_filter_inst_lpf_i_n84, 
      lpf_filter_inst_lpf_i_n83, lpf_filter_inst_lpf_i_n82, 
      lpf_filter_inst_lpf_i_n81, lpf_filter_inst_lpf_i_n80, 
      lpf_filter_inst_lpf_i_n79, lpf_filter_inst_lpf_i_n78, 
      lpf_filter_inst_lpf_i_n77, lpf_filter_inst_lpf_i_n76, 
      lpf_filter_inst_lpf_i_n75, lpf_filter_inst_lpf_i_n74, 
      lpf_filter_inst_lpf_i_n67, lpf_filter_inst_lpf_i_n66, 
      lpf_filter_inst_lpf_i_n65, lpf_filter_inst_lpf_i_n64, 
      lpf_filter_inst_lpf_i_n63, lpf_filter_inst_lpf_i_n62, 
      lpf_filter_inst_lpf_i_n61, lpf_filter_inst_lpf_i_n60, 
      lpf_filter_inst_lpf_i_n59, lpf_filter_inst_lpf_i_n58, 
      lpf_filter_inst_lpf_i_n57, lpf_filter_inst_lpf_i_n56, 
      lpf_filter_inst_lpf_i_n55, lpf_filter_inst_lpf_i_n54, 
      lpf_filter_inst_lpf_i_n53, lpf_filter_inst_lpf_i_n52, 
      lpf_filter_inst_lpf_i_n51, lpf_filter_inst_lpf_i_n50, 
      lpf_filter_inst_lpf_i_n49, lpf_filter_inst_lpf_i_n48, 
      lpf_filter_inst_lpf_i_n47, lpf_filter_inst_lpf_i_n46, 
      lpf_filter_inst_lpf_i_n45, lpf_filter_inst_lpf_i_n44, 
      lpf_filter_inst_lpf_i_n43, lpf_filter_inst_lpf_i_n42, 
      lpf_filter_inst_lpf_i_n41, lpf_filter_inst_lpf_i_n40, 
      lpf_filter_inst_lpf_i_n39, lpf_filter_inst_lpf_i_n38, 
      lpf_filter_inst_lpf_i_n37, lpf_filter_inst_lpf_i_n36, 
      lpf_filter_inst_lpf_i_n35, lpf_filter_inst_lpf_i_n34, 
      lpf_filter_inst_lpf_i_n33, lpf_filter_inst_lpf_i_n32, 
      lpf_filter_inst_lpf_i_n31, lpf_filter_inst_lpf_i_n30, 
      lpf_filter_inst_lpf_i_n29, lpf_filter_inst_lpf_i_n28, 
      lpf_filter_inst_lpf_i_n27, lpf_filter_inst_lpf_i_n26, 
      lpf_filter_inst_lpf_i_n25, lpf_filter_inst_lpf_i_n24, 
      lpf_filter_inst_lpf_i_n23, lpf_filter_inst_lpf_i_n22, 
      lpf_filter_inst_lpf_i_n21, lpf_filter_inst_lpf_i_n20, 
      lpf_filter_inst_lpf_i_n19, lpf_filter_inst_lpf_i_n18, 
      lpf_filter_inst_lpf_i_n17, lpf_filter_inst_lpf_i_n16, 
      lpf_filter_inst_lpf_i_n15, lpf_filter_inst_lpf_i_n14, 
      lpf_filter_inst_lpf_i_n13, lpf_filter_inst_lpf_i_n12, 
      lpf_filter_inst_lpf_i_n11, lpf_filter_inst_lpf_i_n10, 
      lpf_filter_inst_lpf_i_n9, lpf_filter_inst_lpf_i_n8, 
      lpf_filter_inst_lpf_i_n7, lpf_filter_inst_lpf_i_n6, 
      lpf_filter_inst_lpf_i_n5, lpf_filter_inst_lpf_i_n4, 
      lpf_filter_inst_lpf_i_n3, lpf_filter_inst_lpf_i_n2, 
      lpf_filter_inst_lpf_i_n1, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_20_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_19_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_18_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_17_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_16_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_15_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_14_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_13_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_12_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_11_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_10_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_9_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_8_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_7_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_6_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_5_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_4_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_3_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_2_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_11, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_10, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_9, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_8, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_7, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_6, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_5, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_4, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_3, 
      lpf_filter_inst_lpf_i_add_1_root_add_286_carry_2, 
      lpf_filter_inst_lpf_i_sub_280_carry_18_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_17_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_16_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_15_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_14_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_13_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_12_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_11_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_10_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_9_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_8_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_7_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_6_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_5_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_4_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_3_port, 
      lpf_filter_inst_lpf_i_sub_280_carry_2_port, 
      lpf_filter_inst_lpf_i_add_284_carry_13, 
      lpf_filter_inst_lpf_i_add_284_carry_12, 
      lpf_filter_inst_lpf_i_add_284_carry_11, 
      lpf_filter_inst_lpf_i_add_284_carry_10, 
      lpf_filter_inst_lpf_i_add_284_carry_9, 
      lpf_filter_inst_lpf_i_add_284_carry_8, 
      lpf_filter_inst_lpf_i_add_284_carry_7, 
      lpf_filter_inst_lpf_i_add_284_carry_6, 
      lpf_filter_inst_lpf_i_add_284_carry_5, 
      lpf_filter_inst_lpf_i_add_284_carry_4, 
      lpf_filter_inst_lpf_i_add_284_carry_3, lpf_filter_inst_lpf_i_pair3_25_10,
      lpf_filter_inst_lpf_i_pair3_25_11, lpf_filter_inst_lpf_i_pair3_25_12, 
      lpf_filter_inst_lpf_i_pair3_25_2, lpf_filter_inst_lpf_i_pair3_25_3, 
      lpf_filter_inst_lpf_i_pair3_25_4, lpf_filter_inst_lpf_i_pair3_25_5, 
      lpf_filter_inst_lpf_i_pair3_25_6, lpf_filter_inst_lpf_i_pair3_25_7, 
      lpf_filter_inst_lpf_i_pair3_25_8, lpf_filter_inst_lpf_i_pair3_25_9, 
      lpf_filter_inst_lpf_i_pair8_20_0, lpf_filter_inst_lpf_i_pair8_20_10, 
      lpf_filter_inst_lpf_i_pair8_20_11, lpf_filter_inst_lpf_i_pair8_20_12, 
      lpf_filter_inst_lpf_i_pair8_20_1, lpf_filter_inst_lpf_i_pair8_20_2, 
      lpf_filter_inst_lpf_i_pair8_20_3, lpf_filter_inst_lpf_i_pair8_20_4, 
      lpf_filter_inst_lpf_i_pair8_20_5, lpf_filter_inst_lpf_i_pair8_20_6, 
      lpf_filter_inst_lpf_i_pair8_20_7, lpf_filter_inst_lpf_i_pair8_20_8, 
      lpf_filter_inst_lpf_i_pair8_20_9, lpf_filter_inst_lpf_i_pair9_19_0, 
      lpf_filter_inst_lpf_i_pair9_19_10, lpf_filter_inst_lpf_i_pair9_19_11, 
      lpf_filter_inst_lpf_i_pair9_19_12, lpf_filter_inst_lpf_i_pair9_19_1, 
      lpf_filter_inst_lpf_i_pair9_19_2, lpf_filter_inst_lpf_i_pair9_19_3, 
      lpf_filter_inst_lpf_i_pair9_19_4, lpf_filter_inst_lpf_i_pair9_19_5, 
      lpf_filter_inst_lpf_i_pair9_19_6, lpf_filter_inst_lpf_i_pair9_19_7, 
      lpf_filter_inst_lpf_i_pair9_19_8, lpf_filter_inst_lpf_i_pair9_19_9, 
      lpf_filter_inst_lpf_i_p232_2_10, lpf_filter_inst_lpf_i_p232_2_11, 
      lpf_filter_inst_lpf_i_p232_2_12, lpf_filter_inst_lpf_i_p232_2_17, 
      lpf_filter_inst_lpf_i_p232_2_1, lpf_filter_inst_lpf_i_p232_2_2, 
      lpf_filter_inst_lpf_i_p232_2_3, lpf_filter_inst_lpf_i_p232_2_4, 
      lpf_filter_inst_lpf_i_p232_2_5, lpf_filter_inst_lpf_i_p232_2_6, 
      lpf_filter_inst_lpf_i_p232_2_7, lpf_filter_inst_lpf_i_p232_2_8, 
      lpf_filter_inst_lpf_i_p232_2_9, lpf_filter_inst_lpf_i_pair4_24_0, 
      lpf_filter_inst_lpf_i_pair4_24_10, lpf_filter_inst_lpf_i_pair4_24_11, 
      lpf_filter_inst_lpf_i_pair4_24_12, lpf_filter_inst_lpf_i_pair4_24_1, 
      lpf_filter_inst_lpf_i_pair4_24_2, lpf_filter_inst_lpf_i_pair4_24_3, 
      lpf_filter_inst_lpf_i_pair4_24_4, lpf_filter_inst_lpf_i_pair4_24_5, 
      lpf_filter_inst_lpf_i_pair4_24_6, lpf_filter_inst_lpf_i_pair4_24_7, 
      lpf_filter_inst_lpf_i_pair4_24_8, lpf_filter_inst_lpf_i_pair4_24_9, 
      lpf_filter_inst_lpf_i_pair5_23_0, lpf_filter_inst_lpf_i_pair5_23_10, 
      lpf_filter_inst_lpf_i_pair5_23_11, lpf_filter_inst_lpf_i_pair5_23_12, 
      lpf_filter_inst_lpf_i_pair5_23_1, lpf_filter_inst_lpf_i_pair5_23_2, 
      lpf_filter_inst_lpf_i_pair5_23_3, lpf_filter_inst_lpf_i_pair5_23_4, 
      lpf_filter_inst_lpf_i_pair5_23_5, lpf_filter_inst_lpf_i_pair5_23_6, 
      lpf_filter_inst_lpf_i_pair5_23_7, lpf_filter_inst_lpf_i_pair5_23_8, 
      lpf_filter_inst_lpf_i_pair5_23_9, lpf_filter_inst_lpf_i_t4_5_10, 
      lpf_filter_inst_lpf_i_t4_5_11, lpf_filter_inst_lpf_i_t4_5_12, 
      lpf_filter_inst_lpf_i_t4_5_13, lpf_filter_inst_lpf_i_t4_5_2, 
      lpf_filter_inst_lpf_i_t4_5_3, lpf_filter_inst_lpf_i_t4_5_4, 
      lpf_filter_inst_lpf_i_t4_5_5, lpf_filter_inst_lpf_i_t4_5_6, 
      lpf_filter_inst_lpf_i_t4_5_7, lpf_filter_inst_lpf_i_t4_5_8, 
      lpf_filter_inst_lpf_i_t4_5_9, lpf_filter_inst_lpf_i_p206_1_10, 
      lpf_filter_inst_lpf_i_p206_1_11, lpf_filter_inst_lpf_i_p206_1_12, 
      lpf_filter_inst_lpf_i_p206_1_13, lpf_filter_inst_lpf_i_p206_1_14, 
      lpf_filter_inst_lpf_i_p206_1_15, lpf_filter_inst_lpf_i_p206_1_16, 
      lpf_filter_inst_lpf_i_p206_1_17, lpf_filter_inst_lpf_i_p206_1_18, 
      lpf_filter_inst_lpf_i_p206_1_19, lpf_filter_inst_lpf_i_p206_1_3, 
      lpf_filter_inst_lpf_i_p206_1_4, lpf_filter_inst_lpf_i_p206_1_5, 
      lpf_filter_inst_lpf_i_p206_1_6, lpf_filter_inst_lpf_i_p206_1_7, 
      lpf_filter_inst_lpf_i_p206_1_8, lpf_filter_inst_lpf_i_p206_1_9, 
      lpf_filter_inst_lpf_i_pair0_28_0, lpf_filter_inst_lpf_i_pair0_28_10, 
      lpf_filter_inst_lpf_i_pair0_28_11, lpf_filter_inst_lpf_i_pair0_28_12, 
      lpf_filter_inst_lpf_i_pair0_28_1, lpf_filter_inst_lpf_i_pair0_28_2, 
      lpf_filter_inst_lpf_i_pair0_28_3, lpf_filter_inst_lpf_i_pair0_28_4, 
      lpf_filter_inst_lpf_i_pair0_28_5, lpf_filter_inst_lpf_i_pair0_28_6, 
      lpf_filter_inst_lpf_i_pair0_28_7, lpf_filter_inst_lpf_i_pair0_28_8, 
      lpf_filter_inst_lpf_i_pair0_28_9, lpf_filter_inst_lpf_i_t0_1_10, 
      lpf_filter_inst_lpf_i_t0_1_11, lpf_filter_inst_lpf_i_t0_1_12, 
      lpf_filter_inst_lpf_i_t0_1_13, lpf_filter_inst_lpf_i_t0_1_14, 
      lpf_filter_inst_lpf_i_t0_1_1, lpf_filter_inst_lpf_i_t0_1_2, 
      lpf_filter_inst_lpf_i_t0_1_3, lpf_filter_inst_lpf_i_t0_1_4, 
      lpf_filter_inst_lpf_i_t0_1_5, lpf_filter_inst_lpf_i_t0_1_6, 
      lpf_filter_inst_lpf_i_t0_1_7, lpf_filter_inst_lpf_i_t0_1_8, 
      lpf_filter_inst_lpf_i_t0_1_9, lpf_filter_inst_lpf_i_net5306, 
      lpf_filter_inst_lpf_i_t12_13_10, lpf_filter_inst_lpf_i_t12_13_11, 
      lpf_filter_inst_lpf_i_t12_13_12, lpf_filter_inst_lpf_i_t12_13_13, 
      lpf_filter_inst_lpf_i_t12_13_14, lpf_filter_inst_lpf_i_t12_13_15, 
      lpf_filter_inst_lpf_i_t12_13_16, lpf_filter_inst_lpf_i_t12_13_17, 
      lpf_filter_inst_lpf_i_t12_13_18, lpf_filter_inst_lpf_i_t12_13_19, 
      lpf_filter_inst_lpf_i_t12_13_20, lpf_filter_inst_lpf_i_t12_13_21, 
      lpf_filter_inst_lpf_i_t12_13_22, lpf_filter_inst_lpf_i_t12_13_2, 
      lpf_filter_inst_lpf_i_t12_13_3, lpf_filter_inst_lpf_i_t12_13_4, 
      lpf_filter_inst_lpf_i_t12_13_5, lpf_filter_inst_lpf_i_t12_13_6, 
      lpf_filter_inst_lpf_i_t12_13_7, lpf_filter_inst_lpf_i_t12_13_8, 
      lpf_filter_inst_lpf_i_t12_13_9, lpf_filter_inst_lpf_i_n73, 
      lpf_filter_inst_lpf_i_n72, lpf_filter_inst_lpf_i_n71, 
      lpf_filter_inst_lpf_i_n70, lpf_filter_inst_lpf_i_n69, 
      lpf_filter_inst_lpf_i_n68, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_12_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_13_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_14_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_15_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_16_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_17_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_18_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_19_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_20_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_21_port, 
      lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_22_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_3_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_4_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_5_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_6_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_7_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_8_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_9_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_10_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_11_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_12_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_13_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_14_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_15_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_16_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_17_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_18_port, 
      lpf_filter_inst_lpf_i_t4_5_8_9_19_port, 
      lpf_filter_inst_lpf_i_t11_14_0_port, lpf_filter_inst_lpf_i_t11_14_1_port,
      lpf_filter_inst_lpf_i_t11_14_2_port, lpf_filter_inst_lpf_i_t11_14_3_port,
      lpf_filter_inst_lpf_i_t11_14_4_port, lpf_filter_inst_lpf_i_t11_14_5_port,
      lpf_filter_inst_lpf_i_t11_14_6_port, lpf_filter_inst_lpf_i_t11_14_7_port,
      lpf_filter_inst_lpf_i_t11_14_8_port, lpf_filter_inst_lpf_i_t11_14_9_port,
      lpf_filter_inst_lpf_i_t11_14_10_port, 
      lpf_filter_inst_lpf_i_t11_14_11_port, 
      lpf_filter_inst_lpf_i_t11_14_12_port, 
      lpf_filter_inst_lpf_i_t11_14_13_port, 
      lpf_filter_inst_lpf_i_t11_14_14_port, 
      lpf_filter_inst_lpf_i_t11_14_15_port, 
      lpf_filter_inst_lpf_i_t11_14_16_port, 
      lpf_filter_inst_lpf_i_t11_14_17_port, 
      lpf_filter_inst_lpf_i_t11_14_18_port, lpf_filter_inst_lpf_i_p206_3_3_port
      , lpf_filter_inst_lpf_i_p206_3_4_port, 
      lpf_filter_inst_lpf_i_p206_3_5_port, lpf_filter_inst_lpf_i_p206_3_6_port,
      lpf_filter_inst_lpf_i_p206_3_7_port, lpf_filter_inst_lpf_i_p206_3_8_port,
      lpf_filter_inst_lpf_i_p206_3_9_port, lpf_filter_inst_lpf_i_p206_3_10_port
      , lpf_filter_inst_lpf_i_p206_3_11_port, 
      lpf_filter_inst_lpf_i_p206_3_12_port, 
      lpf_filter_inst_lpf_i_p206_3_13_port, 
      lpf_filter_inst_lpf_i_p206_3_14_port, 
      lpf_filter_inst_lpf_i_p206_3_15_port, 
      lpf_filter_inst_lpf_i_p206_3_16_port, 
      lpf_filter_inst_lpf_i_p206_3_17_port, 
      lpf_filter_inst_lpf_i_p206_3_18_port, 
      lpf_filter_inst_lpf_i_p206_3_19_port, 
      lpf_filter_inst_lpf_i_p206_3_20_port, lpf_filter_inst_lpf_i_p206_2_3_port
      , lpf_filter_inst_lpf_i_p206_2_4_port, 
      lpf_filter_inst_lpf_i_p206_2_5_port, lpf_filter_inst_lpf_i_p206_2_6_port,
      lpf_filter_inst_lpf_i_p206_2_7_port, lpf_filter_inst_lpf_i_p206_2_8_port,
      lpf_filter_inst_lpf_i_p206_2_9_port, lpf_filter_inst_lpf_i_p206_2_10_port
      , lpf_filter_inst_lpf_i_p206_2_11_port, 
      lpf_filter_inst_lpf_i_p206_2_12_port, 
      lpf_filter_inst_lpf_i_p206_2_13_port, 
      lpf_filter_inst_lpf_i_p206_2_14_port, 
      lpf_filter_inst_lpf_i_p206_2_15_port, lpf_filter_inst_lpf_i_p141_1_2_port
      , lpf_filter_inst_lpf_i_p141_1_3_port, 
      lpf_filter_inst_lpf_i_p141_1_4_port, lpf_filter_inst_lpf_i_p141_1_5_port,
      lpf_filter_inst_lpf_i_p141_1_6_port, lpf_filter_inst_lpf_i_p141_1_7_port,
      lpf_filter_inst_lpf_i_p141_1_8_port, lpf_filter_inst_lpf_i_p141_1_9_port,
      lpf_filter_inst_lpf_i_p141_1_10_port, 
      lpf_filter_inst_lpf_i_p141_1_11_port, 
      lpf_filter_inst_lpf_i_p141_1_12_port, 
      lpf_filter_inst_lpf_i_p141_1_13_port, 
      lpf_filter_inst_lpf_i_p141_1_14_port, 
      lpf_filter_inst_lpf_i_p141_1_15_port, 
      lpf_filter_inst_lpf_i_p141_1_16_port, 
      lpf_filter_inst_lpf_i_p141_1_17_port, 
      lpf_filter_inst_lpf_i_p141_1_19_port, lpf_filter_inst_lpf_i_t3_7_1_port, 
      lpf_filter_inst_lpf_i_t3_7_2_port, lpf_filter_inst_lpf_i_t3_7_3_port, 
      lpf_filter_inst_lpf_i_t3_7_4_port, lpf_filter_inst_lpf_i_t3_7_5_port, 
      lpf_filter_inst_lpf_i_t3_7_6_port, lpf_filter_inst_lpf_i_t3_7_7_port, 
      lpf_filter_inst_lpf_i_t3_7_8_port, lpf_filter_inst_lpf_i_t3_7_9_port, 
      lpf_filter_inst_lpf_i_t3_7_10_port, lpf_filter_inst_lpf_i_t3_7_11_port, 
      lpf_filter_inst_lpf_i_t3_7_12_port, lpf_filter_inst_lpf_i_t3_7_13_port, 
      lpf_filter_inst_lpf_i_t3_7_14_port, lpf_filter_inst_lpf_i_t3_7_15_port, 
      lpf_filter_inst_lpf_i_t8_9_0_port, lpf_filter_inst_lpf_i_t8_9_1_port, 
      lpf_filter_inst_lpf_i_t8_9_2_port, lpf_filter_inst_lpf_i_t8_9_3_port, 
      lpf_filter_inst_lpf_i_t8_9_4_port, lpf_filter_inst_lpf_i_t8_9_5_port, 
      lpf_filter_inst_lpf_i_t8_9_6_port, lpf_filter_inst_lpf_i_t8_9_7_port, 
      lpf_filter_inst_lpf_i_t8_9_8_port, lpf_filter_inst_lpf_i_t8_9_9_port, 
      lpf_filter_inst_lpf_i_t8_9_10_port, lpf_filter_inst_lpf_i_t8_9_11_port, 
      lpf_filter_inst_lpf_i_t8_9_12_port, lpf_filter_inst_lpf_i_t8_9_13_port, 
      lpf_filter_inst_lpf_i_pair13_15_2_port, 
      lpf_filter_inst_lpf_i_pair13_15_3_port, 
      lpf_filter_inst_lpf_i_pair13_15_4_port, 
      lpf_filter_inst_lpf_i_pair13_15_5_port, 
      lpf_filter_inst_lpf_i_pair13_15_6_port, 
      lpf_filter_inst_lpf_i_pair13_15_7_port, 
      lpf_filter_inst_lpf_i_pair13_15_8_port, 
      lpf_filter_inst_lpf_i_pair13_15_9_port, 
      lpf_filter_inst_lpf_i_pair13_15_10_port, 
      lpf_filter_inst_lpf_i_pair13_15_11_port, 
      lpf_filter_inst_lpf_i_pair12_16_1_port, 
      lpf_filter_inst_lpf_i_pair12_16_2_port, 
      lpf_filter_inst_lpf_i_pair12_16_3_port, 
      lpf_filter_inst_lpf_i_pair12_16_4_port, 
      lpf_filter_inst_lpf_i_pair12_16_5_port, 
      lpf_filter_inst_lpf_i_pair12_16_6_port, 
      lpf_filter_inst_lpf_i_pair12_16_7_port, 
      lpf_filter_inst_lpf_i_pair12_16_8_port, 
      lpf_filter_inst_lpf_i_pair12_16_9_port, 
      lpf_filter_inst_lpf_i_pair12_16_10_port, 
      lpf_filter_inst_lpf_i_pair12_16_11_port, 
      lpf_filter_inst_lpf_i_pair12_16_12_port, 
      lpf_filter_inst_lpf_i_pair11_17_2_port, 
      lpf_filter_inst_lpf_i_pair11_17_3_port, 
      lpf_filter_inst_lpf_i_pair11_17_4_port, 
      lpf_filter_inst_lpf_i_pair11_17_5_port, 
      lpf_filter_inst_lpf_i_pair11_17_6_port, 
      lpf_filter_inst_lpf_i_pair11_17_7_port, 
      lpf_filter_inst_lpf_i_pair11_17_8_port, 
      lpf_filter_inst_lpf_i_pair11_17_9_port, 
      lpf_filter_inst_lpf_i_pair11_17_10_port, 
      lpf_filter_inst_lpf_i_pair11_17_11_port, 
      lpf_filter_inst_lpf_i_pair11_17_12_port, 
      lpf_filter_inst_lpf_i_pair7_21_0_port, 
      lpf_filter_inst_lpf_i_pair7_21_1_port, 
      lpf_filter_inst_lpf_i_pair7_21_2_port, 
      lpf_filter_inst_lpf_i_pair7_21_3_port, 
      lpf_filter_inst_lpf_i_pair7_21_4_port, 
      lpf_filter_inst_lpf_i_pair7_21_5_port, 
      lpf_filter_inst_lpf_i_pair7_21_6_port, 
      lpf_filter_inst_lpf_i_pair7_21_7_port, 
      lpf_filter_inst_lpf_i_pair7_21_8_port, 
      lpf_filter_inst_lpf_i_pair7_21_9_port, 
      lpf_filter_inst_lpf_i_pair7_21_10_port, 
      lpf_filter_inst_lpf_i_pair7_21_11_port, 
      lpf_filter_inst_lpf_i_pair7_21_12_port, 
      lpf_filter_inst_lpf_i_pair1_27_0_port, 
      lpf_filter_inst_lpf_i_pair1_27_1_port, 
      lpf_filter_inst_lpf_i_pair1_27_2_port, 
      lpf_filter_inst_lpf_i_pair1_27_3_port, 
      lpf_filter_inst_lpf_i_pair1_27_4_port, 
      lpf_filter_inst_lpf_i_pair1_27_5_port, 
      lpf_filter_inst_lpf_i_pair1_27_6_port, 
      lpf_filter_inst_lpf_i_pair1_27_7_port, 
      lpf_filter_inst_lpf_i_pair1_27_8_port, 
      lpf_filter_inst_lpf_i_pair1_27_9_port, 
      lpf_filter_inst_lpf_i_pair1_27_10_port, 
      lpf_filter_inst_lpf_i_pair1_27_11_port, 
      lpf_filter_inst_lpf_i_pair1_27_12_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_0_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_1_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_2_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_3_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_4_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_5_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_6_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_7_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_8_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_9_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_10_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_11_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_12_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_13_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_14_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_15_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_16_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_17_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_18_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_19_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_20_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_21_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_22_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_23_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_24_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_25_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_26_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_27_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_28_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_29_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_30_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_31_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_32_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_33_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_34_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_35_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_36_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_37_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_38_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_39_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_40_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_41_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_42_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_43_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_44_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_45_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_46_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_47_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_48_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_49_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_50_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_51_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_52_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_53_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_54_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_55_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_56_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_57_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_58_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_59_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_60_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_61_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_62_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_63_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_64_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_65_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_66_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_67_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_68_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_69_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_70_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_71_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_72_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_73_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_74_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_75_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_76_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_77_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_78_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_79_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_80_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_81_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_82_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_83_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_84_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_85_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_86_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_87_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_88_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_89_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_90_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_91_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_92_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_93_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_94_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_95_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_96_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_97_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_98_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_99_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_100_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_101_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_102_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_103_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_104_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_105_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_106_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_107_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_108_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_109_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_110_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_111_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_112_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_113_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_114_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_115_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_116_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_117_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_118_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_119_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_120_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_121_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_122_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_123_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_124_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_125_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_126_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_127_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_128_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_129_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_130_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_131_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_132_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_133_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_134_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_135_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_136_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_137_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_138_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_139_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_140_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_141_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_142_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_143_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_144_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_145_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_146_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_147_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_148_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_149_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_150_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_151_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_152_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_153_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_154_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_155_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_156_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_157_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_158_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_159_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_160_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_161_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_162_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_163_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_164_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_165_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_166_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_167_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_168_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_169_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_170_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_171_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_172_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_173_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_174_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_175_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_176_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_177_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_178_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_179_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_180_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_181_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_182_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_183_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_184_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_185_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_186_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_187_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_188_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_189_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_190_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_191_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_192_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_193_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_194_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_195_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_196_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_197_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_198_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_199_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_200_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_201_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_202_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_203_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_204_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_205_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_206_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_207_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_208_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_209_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_210_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_211_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_212_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_213_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_214_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_215_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_216_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_217_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_218_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_219_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_220_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_221_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_222_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_223_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_224_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_225_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_226_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_227_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_228_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_229_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_230_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_231_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_232_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_233_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_234_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_235_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_236_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_237_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_238_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_239_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_240_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_241_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_242_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_243_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_244_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_245_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_246_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_247_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_248_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_249_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_250_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_251_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_252_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_253_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_254_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_255_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_256_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_257_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_258_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_259_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_260_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_261_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_262_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_263_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_264_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_265_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_266_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_267_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_268_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_269_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_270_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_271_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_272_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_273_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_274_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_275_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_276_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_277_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_278_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_279_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_280_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_281_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_282_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_283_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_284_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_285_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_286_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_287_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_288_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_289_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_290_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_291_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_292_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_293_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_294_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_295_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_296_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_297_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_298_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_299_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_300_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_301_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_302_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_303_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_304_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_305_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_306_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_307_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_308_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_309_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_310_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_311_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_312_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_313_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_314_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_315_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_316_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_317_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_318_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_319_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_320_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_321_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_322_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_323_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_324_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_325_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_326_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_327_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_328_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_329_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_330_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_331_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_332_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_333_port, 
      lpf_filter_inst_lpf_i_arx_input_reg_334_port, 
      lpf_filter_inst_lpf_i_add_273_n_1308, lpf_filter_inst_lpf_i_add_273_n1, 
      lpf_filter_inst_lpf_i_add_273_carry_2_port, 
      lpf_filter_inst_lpf_i_add_273_carry_3_port, 
      lpf_filter_inst_lpf_i_add_273_carry_4_port, 
      lpf_filter_inst_lpf_i_add_273_carry_5_port, 
      lpf_filter_inst_lpf_i_add_273_carry_6_port, 
      lpf_filter_inst_lpf_i_add_273_carry_7_port, 
      lpf_filter_inst_lpf_i_add_273_carry_8_port, 
      lpf_filter_inst_lpf_i_add_273_carry_9_port, 
      lpf_filter_inst_lpf_i_add_273_carry_10_port, 
      lpf_filter_inst_lpf_i_add_273_carry_11_port, 
      lpf_filter_inst_lpf_i_add_273_carry_12_port, 
      lpf_filter_inst_lpf_i_add_272_n1, 
      lpf_filter_inst_lpf_i_add_272_carry_2_port, 
      lpf_filter_inst_lpf_i_add_272_carry_3_port, 
      lpf_filter_inst_lpf_i_add_272_carry_4_port, 
      lpf_filter_inst_lpf_i_add_272_carry_5_port, 
      lpf_filter_inst_lpf_i_add_272_carry_6_port, 
      lpf_filter_inst_lpf_i_add_272_carry_7_port, 
      lpf_filter_inst_lpf_i_add_272_carry_8_port, 
      lpf_filter_inst_lpf_i_add_272_carry_9_port, 
      lpf_filter_inst_lpf_i_add_272_carry_10_port, 
      lpf_filter_inst_lpf_i_add_272_carry_11_port, 
      lpf_filter_inst_lpf_i_add_272_carry_12_port, 
      lpf_filter_inst_lpf_i_add_271_n_1303, lpf_filter_inst_lpf_i_add_271_n1, 
      lpf_filter_inst_lpf_i_add_271_carry_2_port, 
      lpf_filter_inst_lpf_i_add_271_carry_3_port, 
      lpf_filter_inst_lpf_i_add_271_carry_4_port, 
      lpf_filter_inst_lpf_i_add_271_carry_5_port, 
      lpf_filter_inst_lpf_i_add_271_carry_6_port, 
      lpf_filter_inst_lpf_i_add_271_carry_7_port, 
      lpf_filter_inst_lpf_i_add_271_carry_8_port, 
      lpf_filter_inst_lpf_i_add_271_carry_9_port, 
      lpf_filter_inst_lpf_i_add_271_carry_10_port, 
      lpf_filter_inst_lpf_i_add_271_carry_11_port, 
      lpf_filter_inst_lpf_i_add_271_carry_12_port, 
      lpf_filter_inst_lpf_i_add_268_n1, 
      lpf_filter_inst_lpf_i_add_268_carry_2_port, 
      lpf_filter_inst_lpf_i_add_268_carry_3_port, 
      lpf_filter_inst_lpf_i_add_268_carry_4_port, 
      lpf_filter_inst_lpf_i_add_268_carry_5_port, 
      lpf_filter_inst_lpf_i_add_268_carry_6_port, 
      lpf_filter_inst_lpf_i_add_268_carry_7_port, 
      lpf_filter_inst_lpf_i_add_268_carry_8_port, 
      lpf_filter_inst_lpf_i_add_268_carry_9_port, 
      lpf_filter_inst_lpf_i_add_268_carry_10_port, 
      lpf_filter_inst_lpf_i_add_268_carry_11_port, 
      lpf_filter_inst_lpf_i_add_268_carry_12_port, 
      lpf_filter_inst_lpf_i_add_264_n_1298, lpf_filter_inst_lpf_i_add_264_n1, 
      lpf_filter_inst_lpf_i_add_264_carry_2_port, 
      lpf_filter_inst_lpf_i_add_264_carry_3_port, 
      lpf_filter_inst_lpf_i_add_264_carry_4_port, 
      lpf_filter_inst_lpf_i_add_264_carry_5_port, 
      lpf_filter_inst_lpf_i_add_264_carry_6_port, 
      lpf_filter_inst_lpf_i_add_264_carry_7_port, 
      lpf_filter_inst_lpf_i_add_264_carry_8_port, 
      lpf_filter_inst_lpf_i_add_264_carry_9_port, 
      lpf_filter_inst_lpf_i_add_264_carry_10_port, 
      lpf_filter_inst_lpf_i_add_264_carry_11_port, 
      lpf_filter_inst_lpf_i_add_264_carry_12_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_n1, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_2_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_i_add_5_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_n1, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_i_add_4_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_n_1017, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_n1, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_i_add_7_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_n_1027, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_n1, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_i_add_8_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_n_1036, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_n1, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_i_add_6_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_n_1042, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_n1, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_23_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n_1047, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n16, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n15, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n14, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n13, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n12, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n11, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n10, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n9, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n8, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n7, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n6, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n5, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n4, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n3, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n1, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_23_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_n_1051, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_n1, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_23_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n_1066, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n29, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n28, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n27, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n26, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n25, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n24, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n23, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n22, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n21, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n20, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n19, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n18, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n17, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n16, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n15, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n14, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n13, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n12, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n11, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n10, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n9, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n8, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n7, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n6, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n5, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n4, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n3, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n2, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_23_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_n_1143, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_n1, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_8_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_9_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_10_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_11_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_12_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_13_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_14_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_15_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_16_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_17_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_18_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_285_carry_19_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_n_1254, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_n1, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_2_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_3_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_4_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_5_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_6_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_7_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_8_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_9_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_10_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_11_port, 
      lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_12_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_n_1257, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_n1, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_2_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_3_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_4_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_5_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_6_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_7_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_8_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_9_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_10_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_11_port, 
      lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_12_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_n_1260, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_n1, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_2_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_3_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_4_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_5_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_6_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_7_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_8_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_9_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_10_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_11_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_12_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_13_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n_1265, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n15, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n14, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n13, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n12, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n11, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n10, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n9, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n8, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n7, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n6, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n5, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n4, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n3, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n2, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_n1, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_3_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_4_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_5_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_6_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_7_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_8_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_9_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_10_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_11_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_12_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_13_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_14_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_15_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_16_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_n_1180, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_n1, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_7_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_8_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_9_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_10_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_11_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_12_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_13_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_14_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_15_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_16_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_286_carry_17_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n_1186, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n20, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n19, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n18, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n17, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n16, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n15, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n14, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n13, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n12, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n11, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n10, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n9, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n8, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n7, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n6, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n5, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n4, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n3, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n2, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_n1, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_4_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_5_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_6_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_7_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_8_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_9_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_10_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_11_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_12_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_13_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_14_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_15_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_16_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_17_port, 
      lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_18_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_n_1282, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_n1, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_2_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_3_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_4_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_5_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_6_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_7_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_8_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_9_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_10_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_11_port, 
      lpf_filter_inst_lpf_i_add_1_root_add_277_carry_12_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_n_1285, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_n1, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_2_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_3_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_4_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_5_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_6_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_7_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_8_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_9_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_10_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_11_port, 
      lpf_filter_inst_lpf_i_add_2_root_add_277_carry_12_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_n1, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_2_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_3_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_4_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_5_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_6_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_7_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_8_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_9_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_10_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_11_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_12_port, 
      lpf_filter_inst_lpf_i_add_0_root_add_277_carry_13_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_n_1161, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_n1, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_2_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_3_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_4_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_5_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_6_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_7_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_8_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_9_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_10_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_11_port, 
      lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_12_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n_1166, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n14, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n13, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n12, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n11, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n10, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n9, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n8, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n7, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n6, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n5, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n4, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n3, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n2, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_n1, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_3_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_4_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_5_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_6_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_7_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_8_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_9_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_10_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_11_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_12_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_13_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_14_port, 
      lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_15_port, 
      lpf_filter_inst_lpf_q_n_1371, lpf_filter_inst_lpf_q_n_1370, 
      lpf_filter_inst_lpf_q_n_1369, lpf_filter_inst_lpf_q_n_1368, 
      lpf_filter_inst_lpf_q_n_1367, lpf_filter_inst_lpf_q_n_1366, 
      lpf_filter_inst_lpf_q_n_1365, lpf_filter_inst_lpf_q_n_1364, 
      lpf_filter_inst_lpf_q_n_1363, lpf_filter_inst_lpf_q_n_1362, 
      lpf_filter_inst_lpf_q_n_1361, lpf_filter_inst_lpf_q_n_1360, 
      lpf_filter_inst_lpf_q_n_1359, lpf_filter_inst_lpf_q_n_1358, 
      lpf_filter_inst_lpf_q_n_1357, lpf_filter_inst_lpf_q_n_1356, 
      lpf_filter_inst_lpf_q_n_1355, lpf_filter_inst_lpf_q_n_1354, 
      lpf_filter_inst_lpf_q_n_1353, lpf_filter_inst_lpf_q_n_1352, 
      lpf_filter_inst_lpf_q_n_1351, lpf_filter_inst_lpf_q_n_1350, 
      lpf_filter_inst_lpf_q_n_1349, lpf_filter_inst_lpf_q_n_1348, 
      lpf_filter_inst_lpf_q_n_1347, lpf_filter_inst_lpf_q_n_1346, 
      lpf_filter_inst_lpf_q_n_1345, lpf_filter_inst_lpf_q_n_1344, 
      lpf_filter_inst_lpf_q_n_1343, lpf_filter_inst_lpf_q_n_1342, 
      lpf_filter_inst_lpf_q_n_1341, lpf_filter_inst_lpf_q_n_1340, 
      lpf_filter_inst_lpf_q_n_1339, lpf_filter_inst_lpf_q_n_1338, 
      lpf_filter_inst_lpf_q_n_1337, lpf_filter_inst_lpf_q_n_1336, 
      lpf_filter_inst_lpf_q_n_1335, lpf_filter_inst_lpf_q_n_1334, 
      lpf_filter_inst_lpf_q_n_1333, lpf_filter_inst_lpf_q_n_1332, 
      lpf_filter_inst_lpf_q_n_1331, lpf_filter_inst_lpf_q_n_1330, 
      lpf_filter_inst_lpf_q_n_1329, lpf_filter_inst_lpf_q_n_1328, 
      lpf_filter_inst_lpf_q_n_1327, lpf_filter_inst_lpf_q_n_1326, 
      lpf_filter_inst_lpf_q_n_1325, lpf_filter_inst_lpf_q_n_1324, 
      lpf_filter_inst_lpf_q_n_1323, lpf_filter_inst_lpf_q_n_1322, 
      lpf_filter_inst_lpf_q_n200, lpf_filter_inst_lpf_q_n199, 
      lpf_filter_inst_lpf_q_n198, lpf_filter_inst_lpf_q_n197, 
      lpf_filter_inst_lpf_q_n196, lpf_filter_inst_lpf_q_n195, 
      lpf_filter_inst_lpf_q_n194, lpf_filter_inst_lpf_q_n193, 
      lpf_filter_inst_lpf_q_n192, lpf_filter_inst_lpf_q_n191, 
      lpf_filter_inst_lpf_q_n190, lpf_filter_inst_lpf_q_n189, 
      lpf_filter_inst_lpf_q_n188, lpf_filter_inst_lpf_q_n187, 
      lpf_filter_inst_lpf_q_n186, lpf_filter_inst_lpf_q_n185, 
      lpf_filter_inst_lpf_q_n184, lpf_filter_inst_lpf_q_n183, 
      lpf_filter_inst_lpf_q_n182, lpf_filter_inst_lpf_q_n181, 
      lpf_filter_inst_lpf_q_n180, lpf_filter_inst_lpf_q_n179, 
      lpf_filter_inst_lpf_q_n178, lpf_filter_inst_lpf_q_n177, 
      lpf_filter_inst_lpf_q_n176, lpf_filter_inst_lpf_q_n175, 
      lpf_filter_inst_lpf_q_n174, lpf_filter_inst_lpf_q_n173, 
      lpf_filter_inst_lpf_q_n172, lpf_filter_inst_lpf_q_n171, 
      lpf_filter_inst_lpf_q_n170, lpf_filter_inst_lpf_q_n169, 
      lpf_filter_inst_lpf_q_n168, lpf_filter_inst_lpf_q_n167, 
      lpf_filter_inst_lpf_q_n166, lpf_filter_inst_lpf_q_n165, 
      lpf_filter_inst_lpf_q_n164, lpf_filter_inst_lpf_q_n163, 
      lpf_filter_inst_lpf_q_n162, lpf_filter_inst_lpf_q_n161, 
      lpf_filter_inst_lpf_q_n160, lpf_filter_inst_lpf_q_n159, 
      lpf_filter_inst_lpf_q_n157, lpf_filter_inst_lpf_q_n156, 
      lpf_filter_inst_lpf_q_n155, lpf_filter_inst_lpf_q_n154, 
      lpf_filter_inst_lpf_q_n153, lpf_filter_inst_lpf_q_n152, 
      lpf_filter_inst_lpf_q_n151, lpf_filter_inst_lpf_q_n150, 
      lpf_filter_inst_lpf_q_n149, lpf_filter_inst_lpf_q_n148, 
      lpf_filter_inst_lpf_q_n147, lpf_filter_inst_lpf_q_n146, 
      lpf_filter_inst_lpf_q_n145, lpf_filter_inst_lpf_q_n144, 
      lpf_filter_inst_lpf_q_n143, lpf_filter_inst_lpf_q_n142, 
      lpf_filter_inst_lpf_q_n141, lpf_filter_inst_lpf_q_n140, 
      lpf_filter_inst_lpf_q_n139, lpf_filter_inst_lpf_q_n138, 
      lpf_filter_inst_lpf_q_n137, lpf_filter_inst_lpf_q_n136, 
      lpf_filter_inst_lpf_q_n135, lpf_filter_inst_lpf_q_n134, 
      lpf_filter_inst_lpf_q_n133, lpf_filter_inst_lpf_q_n132, 
      lpf_filter_inst_lpf_q_n131, lpf_filter_inst_lpf_q_n130, 
      lpf_filter_inst_lpf_q_n129, lpf_filter_inst_lpf_q_n128, 
      lpf_filter_inst_lpf_q_n127, lpf_filter_inst_lpf_q_n126, 
      lpf_filter_inst_lpf_q_n125, lpf_filter_inst_lpf_q_n124, 
      lpf_filter_inst_lpf_q_n123, lpf_filter_inst_lpf_q_n122, 
      lpf_filter_inst_lpf_q_n121, lpf_filter_inst_lpf_q_n120, 
      lpf_filter_inst_lpf_q_n119, lpf_filter_inst_lpf_q_n118, 
      lpf_filter_inst_lpf_q_n117, lpf_filter_inst_lpf_q_n116, 
      lpf_filter_inst_lpf_q_n115, lpf_filter_inst_lpf_q_n114, 
      lpf_filter_inst_lpf_q_n113, lpf_filter_inst_lpf_q_n112, 
      lpf_filter_inst_lpf_q_n111, lpf_filter_inst_lpf_q_n110, 
      lpf_filter_inst_lpf_q_n109, lpf_filter_inst_lpf_q_n108, 
      lpf_filter_inst_lpf_q_n107, lpf_filter_inst_lpf_q_n106, 
      lpf_filter_inst_lpf_q_n105, lpf_filter_inst_lpf_q_n104, 
      lpf_filter_inst_lpf_q_n103, lpf_filter_inst_lpf_q_n102, 
      lpf_filter_inst_lpf_q_n101, lpf_filter_inst_lpf_q_n100, 
      lpf_filter_inst_lpf_q_n99, lpf_filter_inst_lpf_q_n98, 
      lpf_filter_inst_lpf_q_n97, lpf_filter_inst_lpf_q_n96, 
      lpf_filter_inst_lpf_q_n95, lpf_filter_inst_lpf_q_n94, 
      lpf_filter_inst_lpf_q_n92, lpf_filter_inst_lpf_q_n91, 
      lpf_filter_inst_lpf_q_n90, lpf_filter_inst_lpf_q_n89, 
      lpf_filter_inst_lpf_q_n88, lpf_filter_inst_lpf_q_n87, 
      lpf_filter_inst_lpf_q_n86, lpf_filter_inst_lpf_q_n85, 
      lpf_filter_inst_lpf_q_n84, lpf_filter_inst_lpf_q_n83, 
      lpf_filter_inst_lpf_q_n82, lpf_filter_inst_lpf_q_n81, 
      lpf_filter_inst_lpf_q_n80, lpf_filter_inst_lpf_q_n79, 
      lpf_filter_inst_lpf_q_n78, lpf_filter_inst_lpf_q_n77, 
      lpf_filter_inst_lpf_q_n76, lpf_filter_inst_lpf_q_n75, 
      lpf_filter_inst_lpf_q_n74, lpf_filter_inst_lpf_q_n67, 
      lpf_filter_inst_lpf_q_n66, lpf_filter_inst_lpf_q_n65, 
      lpf_filter_inst_lpf_q_n64, lpf_filter_inst_lpf_q_n63, 
      lpf_filter_inst_lpf_q_n62, lpf_filter_inst_lpf_q_n61, 
      lpf_filter_inst_lpf_q_n60, lpf_filter_inst_lpf_q_n59, 
      lpf_filter_inst_lpf_q_n58, lpf_filter_inst_lpf_q_n57, 
      lpf_filter_inst_lpf_q_n56, lpf_filter_inst_lpf_q_n55, 
      lpf_filter_inst_lpf_q_n54, lpf_filter_inst_lpf_q_n53, 
      lpf_filter_inst_lpf_q_n52, lpf_filter_inst_lpf_q_n51, 
      lpf_filter_inst_lpf_q_n50, lpf_filter_inst_lpf_q_n49, 
      lpf_filter_inst_lpf_q_n48, lpf_filter_inst_lpf_q_n47, 
      lpf_filter_inst_lpf_q_n46, lpf_filter_inst_lpf_q_n45, 
      lpf_filter_inst_lpf_q_n44, lpf_filter_inst_lpf_q_n43, 
      lpf_filter_inst_lpf_q_n42, lpf_filter_inst_lpf_q_n41, 
      lpf_filter_inst_lpf_q_n40, lpf_filter_inst_lpf_q_n39, 
      lpf_filter_inst_lpf_q_n38, lpf_filter_inst_lpf_q_n37, 
      lpf_filter_inst_lpf_q_n36, lpf_filter_inst_lpf_q_n35, 
      lpf_filter_inst_lpf_q_n34, lpf_filter_inst_lpf_q_n33, 
      lpf_filter_inst_lpf_q_n32, lpf_filter_inst_lpf_q_n31, 
      lpf_filter_inst_lpf_q_n30, lpf_filter_inst_lpf_q_n29, 
      lpf_filter_inst_lpf_q_n28, lpf_filter_inst_lpf_q_n27, 
      lpf_filter_inst_lpf_q_n26, lpf_filter_inst_lpf_q_n25, 
      lpf_filter_inst_lpf_q_n24, lpf_filter_inst_lpf_q_n23, 
      lpf_filter_inst_lpf_q_n22, lpf_filter_inst_lpf_q_n21, 
      lpf_filter_inst_lpf_q_n20, lpf_filter_inst_lpf_q_n19, 
      lpf_filter_inst_lpf_q_n18, lpf_filter_inst_lpf_q_n17, 
      lpf_filter_inst_lpf_q_n16, lpf_filter_inst_lpf_q_n15, 
      lpf_filter_inst_lpf_q_n14, lpf_filter_inst_lpf_q_n13, 
      lpf_filter_inst_lpf_q_n12, lpf_filter_inst_lpf_q_n11, 
      lpf_filter_inst_lpf_q_n10, lpf_filter_inst_lpf_q_n9, 
      lpf_filter_inst_lpf_q_n8, lpf_filter_inst_lpf_q_n7, 
      lpf_filter_inst_lpf_q_n6, lpf_filter_inst_lpf_q_n5, 
      lpf_filter_inst_lpf_q_n4, lpf_filter_inst_lpf_q_n3, 
      lpf_filter_inst_lpf_q_n2, lpf_filter_inst_lpf_q_n1, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_20_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_19_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_18_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_17_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_16_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_15_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_14_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_13_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_12_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_11_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_10_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_9_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_8_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_7_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_6_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_5_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_4_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_3_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_2_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_11, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_10, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_9, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_8, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_7, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_6, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_5, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_4, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_3, 
      lpf_filter_inst_lpf_q_add_1_root_add_286_carry_2, 
      lpf_filter_inst_lpf_q_sub_280_carry_18_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_17_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_16_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_15_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_14_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_13_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_12_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_11_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_10_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_9_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_8_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_7_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_6_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_5_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_4_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_3_port, 
      lpf_filter_inst_lpf_q_sub_280_carry_2_port, 
      lpf_filter_inst_lpf_q_add_284_carry_13, 
      lpf_filter_inst_lpf_q_add_284_carry_12, 
      lpf_filter_inst_lpf_q_add_284_carry_11, 
      lpf_filter_inst_lpf_q_add_284_carry_10, 
      lpf_filter_inst_lpf_q_add_284_carry_9, 
      lpf_filter_inst_lpf_q_add_284_carry_8, 
      lpf_filter_inst_lpf_q_add_284_carry_7, 
      lpf_filter_inst_lpf_q_add_284_carry_6, 
      lpf_filter_inst_lpf_q_add_284_carry_5, 
      lpf_filter_inst_lpf_q_add_284_carry_4, 
      lpf_filter_inst_lpf_q_add_284_carry_3, lpf_filter_inst_lpf_q_pair3_25_10,
      lpf_filter_inst_lpf_q_pair3_25_11, lpf_filter_inst_lpf_q_pair3_25_12, 
      lpf_filter_inst_lpf_q_pair3_25_2, lpf_filter_inst_lpf_q_pair3_25_3, 
      lpf_filter_inst_lpf_q_pair3_25_4, lpf_filter_inst_lpf_q_pair3_25_5, 
      lpf_filter_inst_lpf_q_pair3_25_6, lpf_filter_inst_lpf_q_pair3_25_7, 
      lpf_filter_inst_lpf_q_pair3_25_8, lpf_filter_inst_lpf_q_pair3_25_9, 
      lpf_filter_inst_lpf_q_pair8_20_0, lpf_filter_inst_lpf_q_pair8_20_10, 
      lpf_filter_inst_lpf_q_pair8_20_11, lpf_filter_inst_lpf_q_pair8_20_12, 
      lpf_filter_inst_lpf_q_pair8_20_1, lpf_filter_inst_lpf_q_pair8_20_2, 
      lpf_filter_inst_lpf_q_pair8_20_3, lpf_filter_inst_lpf_q_pair8_20_4, 
      lpf_filter_inst_lpf_q_pair8_20_5, lpf_filter_inst_lpf_q_pair8_20_6, 
      lpf_filter_inst_lpf_q_pair8_20_7, lpf_filter_inst_lpf_q_pair8_20_8, 
      lpf_filter_inst_lpf_q_pair8_20_9, lpf_filter_inst_lpf_q_pair9_19_0, 
      lpf_filter_inst_lpf_q_pair9_19_10, lpf_filter_inst_lpf_q_pair9_19_11, 
      lpf_filter_inst_lpf_q_pair9_19_12, lpf_filter_inst_lpf_q_pair9_19_1, 
      lpf_filter_inst_lpf_q_pair9_19_2, lpf_filter_inst_lpf_q_pair9_19_3, 
      lpf_filter_inst_lpf_q_pair9_19_4, lpf_filter_inst_lpf_q_pair9_19_5, 
      lpf_filter_inst_lpf_q_pair9_19_6, lpf_filter_inst_lpf_q_pair9_19_7, 
      lpf_filter_inst_lpf_q_pair9_19_8, lpf_filter_inst_lpf_q_pair9_19_9, 
      lpf_filter_inst_lpf_q_p232_2_10, lpf_filter_inst_lpf_q_p232_2_11, 
      lpf_filter_inst_lpf_q_p232_2_12, lpf_filter_inst_lpf_q_p232_2_17, 
      lpf_filter_inst_lpf_q_p232_2_1, lpf_filter_inst_lpf_q_p232_2_2, 
      lpf_filter_inst_lpf_q_p232_2_3, lpf_filter_inst_lpf_q_p232_2_4, 
      lpf_filter_inst_lpf_q_p232_2_5, lpf_filter_inst_lpf_q_p232_2_6, 
      lpf_filter_inst_lpf_q_p232_2_7, lpf_filter_inst_lpf_q_p232_2_8, 
      lpf_filter_inst_lpf_q_p232_2_9, lpf_filter_inst_lpf_q_pair4_24_0, 
      lpf_filter_inst_lpf_q_pair4_24_10, lpf_filter_inst_lpf_q_pair4_24_11, 
      lpf_filter_inst_lpf_q_pair4_24_12, lpf_filter_inst_lpf_q_pair4_24_1, 
      lpf_filter_inst_lpf_q_pair4_24_2, lpf_filter_inst_lpf_q_pair4_24_3, 
      lpf_filter_inst_lpf_q_pair4_24_4, lpf_filter_inst_lpf_q_pair4_24_5, 
      lpf_filter_inst_lpf_q_pair4_24_6, lpf_filter_inst_lpf_q_pair4_24_7, 
      lpf_filter_inst_lpf_q_pair4_24_8, lpf_filter_inst_lpf_q_pair4_24_9, 
      lpf_filter_inst_lpf_q_pair5_23_0, lpf_filter_inst_lpf_q_pair5_23_10, 
      lpf_filter_inst_lpf_q_pair5_23_11, lpf_filter_inst_lpf_q_pair5_23_12, 
      lpf_filter_inst_lpf_q_pair5_23_1, lpf_filter_inst_lpf_q_pair5_23_2, 
      lpf_filter_inst_lpf_q_pair5_23_3, lpf_filter_inst_lpf_q_pair5_23_4, 
      lpf_filter_inst_lpf_q_pair5_23_5, lpf_filter_inst_lpf_q_pair5_23_6, 
      lpf_filter_inst_lpf_q_pair5_23_7, lpf_filter_inst_lpf_q_pair5_23_8, 
      lpf_filter_inst_lpf_q_pair5_23_9, lpf_filter_inst_lpf_q_t4_5_10, 
      lpf_filter_inst_lpf_q_t4_5_11, lpf_filter_inst_lpf_q_t4_5_12, 
      lpf_filter_inst_lpf_q_t4_5_13, lpf_filter_inst_lpf_q_t4_5_2, 
      lpf_filter_inst_lpf_q_t4_5_3, lpf_filter_inst_lpf_q_t4_5_4, 
      lpf_filter_inst_lpf_q_t4_5_5, lpf_filter_inst_lpf_q_t4_5_6, 
      lpf_filter_inst_lpf_q_t4_5_7, lpf_filter_inst_lpf_q_t4_5_8, 
      lpf_filter_inst_lpf_q_t4_5_9, lpf_filter_inst_lpf_q_p206_1_10, 
      lpf_filter_inst_lpf_q_p206_1_11, lpf_filter_inst_lpf_q_p206_1_12, 
      lpf_filter_inst_lpf_q_p206_1_13, lpf_filter_inst_lpf_q_p206_1_14, 
      lpf_filter_inst_lpf_q_p206_1_15, lpf_filter_inst_lpf_q_p206_1_16, 
      lpf_filter_inst_lpf_q_p206_1_17, lpf_filter_inst_lpf_q_p206_1_18, 
      lpf_filter_inst_lpf_q_p206_1_19, lpf_filter_inst_lpf_q_p206_1_3, 
      lpf_filter_inst_lpf_q_p206_1_4, lpf_filter_inst_lpf_q_p206_1_5, 
      lpf_filter_inst_lpf_q_p206_1_6, lpf_filter_inst_lpf_q_p206_1_7, 
      lpf_filter_inst_lpf_q_p206_1_8, lpf_filter_inst_lpf_q_p206_1_9, 
      lpf_filter_inst_lpf_q_pair0_28_0, lpf_filter_inst_lpf_q_pair0_28_10, 
      lpf_filter_inst_lpf_q_pair0_28_11, lpf_filter_inst_lpf_q_pair0_28_12, 
      lpf_filter_inst_lpf_q_pair0_28_1, lpf_filter_inst_lpf_q_pair0_28_2, 
      lpf_filter_inst_lpf_q_pair0_28_3, lpf_filter_inst_lpf_q_pair0_28_4, 
      lpf_filter_inst_lpf_q_pair0_28_5, lpf_filter_inst_lpf_q_pair0_28_6, 
      lpf_filter_inst_lpf_q_pair0_28_7, lpf_filter_inst_lpf_q_pair0_28_8, 
      lpf_filter_inst_lpf_q_pair0_28_9, lpf_filter_inst_lpf_q_t0_1_10, 
      lpf_filter_inst_lpf_q_t0_1_11, lpf_filter_inst_lpf_q_t0_1_12, 
      lpf_filter_inst_lpf_q_t0_1_13, lpf_filter_inst_lpf_q_t0_1_14, 
      lpf_filter_inst_lpf_q_t0_1_1, lpf_filter_inst_lpf_q_t0_1_2, 
      lpf_filter_inst_lpf_q_t0_1_3, lpf_filter_inst_lpf_q_t0_1_4, 
      lpf_filter_inst_lpf_q_t0_1_5, lpf_filter_inst_lpf_q_t0_1_6, 
      lpf_filter_inst_lpf_q_t0_1_7, lpf_filter_inst_lpf_q_t0_1_8, 
      lpf_filter_inst_lpf_q_t0_1_9, lpf_filter_inst_lpf_q_net5308, 
      lpf_filter_inst_lpf_q_t12_13_10, lpf_filter_inst_lpf_q_t12_13_11, 
      lpf_filter_inst_lpf_q_t12_13_12, lpf_filter_inst_lpf_q_t12_13_13, 
      lpf_filter_inst_lpf_q_t12_13_14, lpf_filter_inst_lpf_q_t12_13_15, 
      lpf_filter_inst_lpf_q_t12_13_16, lpf_filter_inst_lpf_q_t12_13_17, 
      lpf_filter_inst_lpf_q_t12_13_18, lpf_filter_inst_lpf_q_t12_13_19, 
      lpf_filter_inst_lpf_q_t12_13_20, lpf_filter_inst_lpf_q_t12_13_21, 
      lpf_filter_inst_lpf_q_t12_13_22, lpf_filter_inst_lpf_q_t12_13_2, 
      lpf_filter_inst_lpf_q_t12_13_3, lpf_filter_inst_lpf_q_t12_13_4, 
      lpf_filter_inst_lpf_q_t12_13_5, lpf_filter_inst_lpf_q_t12_13_6, 
      lpf_filter_inst_lpf_q_t12_13_7, lpf_filter_inst_lpf_q_t12_13_8, 
      lpf_filter_inst_lpf_q_t12_13_9, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_12_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_13_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_14_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_15_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_16_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_17_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_18_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_19_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_20_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_21_port, 
      lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_22_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_3_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_4_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_5_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_6_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_7_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_8_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_9_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_10_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_11_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_12_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_13_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_14_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_15_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_16_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_17_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_18_port, 
      lpf_filter_inst_lpf_q_t4_5_8_9_19_port, 
      lpf_filter_inst_lpf_q_t11_14_0_port, lpf_filter_inst_lpf_q_t11_14_1_port,
      lpf_filter_inst_lpf_q_t11_14_2_port, lpf_filter_inst_lpf_q_t11_14_3_port,
      lpf_filter_inst_lpf_q_t11_14_4_port, lpf_filter_inst_lpf_q_t11_14_5_port,
      lpf_filter_inst_lpf_q_t11_14_6_port, lpf_filter_inst_lpf_q_t11_14_7_port,
      lpf_filter_inst_lpf_q_t11_14_8_port, lpf_filter_inst_lpf_q_t11_14_9_port,
      lpf_filter_inst_lpf_q_t11_14_10_port, 
      lpf_filter_inst_lpf_q_t11_14_11_port, 
      lpf_filter_inst_lpf_q_t11_14_12_port, 
      lpf_filter_inst_lpf_q_t11_14_13_port, 
      lpf_filter_inst_lpf_q_t11_14_14_port, 
      lpf_filter_inst_lpf_q_t11_14_15_port, 
      lpf_filter_inst_lpf_q_t11_14_16_port, 
      lpf_filter_inst_lpf_q_t11_14_17_port, 
      lpf_filter_inst_lpf_q_t11_14_18_port, lpf_filter_inst_lpf_q_p206_3_3_port
      , lpf_filter_inst_lpf_q_p206_3_4_port, 
      lpf_filter_inst_lpf_q_p206_3_5_port, lpf_filter_inst_lpf_q_p206_3_6_port,
      lpf_filter_inst_lpf_q_p206_3_7_port, lpf_filter_inst_lpf_q_p206_3_8_port,
      lpf_filter_inst_lpf_q_p206_3_9_port, lpf_filter_inst_lpf_q_p206_3_10_port
      , lpf_filter_inst_lpf_q_p206_3_11_port, 
      lpf_filter_inst_lpf_q_p206_3_12_port, 
      lpf_filter_inst_lpf_q_p206_3_13_port, 
      lpf_filter_inst_lpf_q_p206_3_14_port, 
      lpf_filter_inst_lpf_q_p206_3_15_port, 
      lpf_filter_inst_lpf_q_p206_3_16_port, 
      lpf_filter_inst_lpf_q_p206_3_17_port, 
      lpf_filter_inst_lpf_q_p206_3_18_port, 
      lpf_filter_inst_lpf_q_p206_3_19_port, 
      lpf_filter_inst_lpf_q_p206_3_20_port, lpf_filter_inst_lpf_q_p206_2_3_port
      , lpf_filter_inst_lpf_q_p206_2_4_port, 
      lpf_filter_inst_lpf_q_p206_2_5_port, lpf_filter_inst_lpf_q_p206_2_6_port,
      lpf_filter_inst_lpf_q_p206_2_7_port, lpf_filter_inst_lpf_q_p206_2_8_port,
      lpf_filter_inst_lpf_q_p206_2_9_port, lpf_filter_inst_lpf_q_p206_2_10_port
      , lpf_filter_inst_lpf_q_p206_2_11_port, 
      lpf_filter_inst_lpf_q_p206_2_12_port, 
      lpf_filter_inst_lpf_q_p206_2_13_port, 
      lpf_filter_inst_lpf_q_p206_2_14_port, 
      lpf_filter_inst_lpf_q_p206_2_15_port, lpf_filter_inst_lpf_q_p141_1_2_port
      , lpf_filter_inst_lpf_q_p141_1_3_port, 
      lpf_filter_inst_lpf_q_p141_1_4_port, lpf_filter_inst_lpf_q_p141_1_5_port,
      lpf_filter_inst_lpf_q_p141_1_6_port, lpf_filter_inst_lpf_q_p141_1_7_port,
      lpf_filter_inst_lpf_q_p141_1_8_port, lpf_filter_inst_lpf_q_p141_1_9_port,
      lpf_filter_inst_lpf_q_p141_1_10_port, 
      lpf_filter_inst_lpf_q_p141_1_11_port, 
      lpf_filter_inst_lpf_q_p141_1_12_port, 
      lpf_filter_inst_lpf_q_p141_1_13_port, 
      lpf_filter_inst_lpf_q_p141_1_14_port, 
      lpf_filter_inst_lpf_q_p141_1_15_port, 
      lpf_filter_inst_lpf_q_p141_1_16_port, 
      lpf_filter_inst_lpf_q_p141_1_17_port, 
      lpf_filter_inst_lpf_q_p141_1_19_port, lpf_filter_inst_lpf_q_t3_7_1_port, 
      lpf_filter_inst_lpf_q_t3_7_2_port, lpf_filter_inst_lpf_q_t3_7_3_port, 
      lpf_filter_inst_lpf_q_t3_7_4_port, lpf_filter_inst_lpf_q_t3_7_5_port, 
      lpf_filter_inst_lpf_q_t3_7_6_port, lpf_filter_inst_lpf_q_t3_7_7_port, 
      lpf_filter_inst_lpf_q_t3_7_8_port, lpf_filter_inst_lpf_q_t3_7_9_port, 
      lpf_filter_inst_lpf_q_t3_7_10_port, lpf_filter_inst_lpf_q_t3_7_11_port, 
      lpf_filter_inst_lpf_q_t3_7_12_port, lpf_filter_inst_lpf_q_t3_7_13_port, 
      lpf_filter_inst_lpf_q_t3_7_14_port, lpf_filter_inst_lpf_q_t3_7_15_port, 
      lpf_filter_inst_lpf_q_t8_9_0_port, lpf_filter_inst_lpf_q_t8_9_1_port, 
      lpf_filter_inst_lpf_q_t8_9_2_port, lpf_filter_inst_lpf_q_t8_9_3_port, 
      lpf_filter_inst_lpf_q_t8_9_4_port, lpf_filter_inst_lpf_q_t8_9_5_port, 
      lpf_filter_inst_lpf_q_t8_9_6_port, lpf_filter_inst_lpf_q_t8_9_7_port, 
      lpf_filter_inst_lpf_q_t8_9_8_port, lpf_filter_inst_lpf_q_t8_9_9_port, 
      lpf_filter_inst_lpf_q_t8_9_10_port, lpf_filter_inst_lpf_q_t8_9_11_port, 
      lpf_filter_inst_lpf_q_t8_9_12_port, lpf_filter_inst_lpf_q_t8_9_13_port, 
      lpf_filter_inst_lpf_q_pair13_15_2_port, 
      lpf_filter_inst_lpf_q_pair13_15_3_port, 
      lpf_filter_inst_lpf_q_pair13_15_4_port, 
      lpf_filter_inst_lpf_q_pair13_15_5_port, 
      lpf_filter_inst_lpf_q_pair13_15_6_port, 
      lpf_filter_inst_lpf_q_pair13_15_7_port, 
      lpf_filter_inst_lpf_q_pair13_15_8_port, 
      lpf_filter_inst_lpf_q_pair13_15_9_port, 
      lpf_filter_inst_lpf_q_pair13_15_10_port, 
      lpf_filter_inst_lpf_q_pair13_15_11_port, 
      lpf_filter_inst_lpf_q_pair12_16_1_port, 
      lpf_filter_inst_lpf_q_pair12_16_2_port, 
      lpf_filter_inst_lpf_q_pair12_16_3_port, 
      lpf_filter_inst_lpf_q_pair12_16_4_port, 
      lpf_filter_inst_lpf_q_pair12_16_5_port, 
      lpf_filter_inst_lpf_q_pair12_16_6_port, 
      lpf_filter_inst_lpf_q_pair12_16_7_port, 
      lpf_filter_inst_lpf_q_pair12_16_8_port, 
      lpf_filter_inst_lpf_q_pair12_16_9_port, 
      lpf_filter_inst_lpf_q_pair12_16_10_port, 
      lpf_filter_inst_lpf_q_pair12_16_11_port, 
      lpf_filter_inst_lpf_q_pair12_16_12_port, 
      lpf_filter_inst_lpf_q_pair11_17_2_port, 
      lpf_filter_inst_lpf_q_pair11_17_3_port, 
      lpf_filter_inst_lpf_q_pair11_17_4_port, 
      lpf_filter_inst_lpf_q_pair11_17_5_port, 
      lpf_filter_inst_lpf_q_pair11_17_6_port, 
      lpf_filter_inst_lpf_q_pair11_17_7_port, 
      lpf_filter_inst_lpf_q_pair11_17_8_port, 
      lpf_filter_inst_lpf_q_pair11_17_9_port, 
      lpf_filter_inst_lpf_q_pair11_17_10_port, 
      lpf_filter_inst_lpf_q_pair11_17_11_port, 
      lpf_filter_inst_lpf_q_pair11_17_12_port, 
      lpf_filter_inst_lpf_q_pair7_21_0_port, 
      lpf_filter_inst_lpf_q_pair7_21_1_port, 
      lpf_filter_inst_lpf_q_pair7_21_2_port, 
      lpf_filter_inst_lpf_q_pair7_21_3_port, 
      lpf_filter_inst_lpf_q_pair7_21_4_port, 
      lpf_filter_inst_lpf_q_pair7_21_5_port, 
      lpf_filter_inst_lpf_q_pair7_21_6_port, 
      lpf_filter_inst_lpf_q_pair7_21_7_port, 
      lpf_filter_inst_lpf_q_pair7_21_8_port, 
      lpf_filter_inst_lpf_q_pair7_21_9_port, 
      lpf_filter_inst_lpf_q_pair7_21_10_port, 
      lpf_filter_inst_lpf_q_pair7_21_11_port, 
      lpf_filter_inst_lpf_q_pair7_21_12_port, 
      lpf_filter_inst_lpf_q_pair1_27_0_port, 
      lpf_filter_inst_lpf_q_pair1_27_1_port, 
      lpf_filter_inst_lpf_q_pair1_27_2_port, 
      lpf_filter_inst_lpf_q_pair1_27_3_port, 
      lpf_filter_inst_lpf_q_pair1_27_4_port, 
      lpf_filter_inst_lpf_q_pair1_27_5_port, 
      lpf_filter_inst_lpf_q_pair1_27_6_port, 
      lpf_filter_inst_lpf_q_pair1_27_7_port, 
      lpf_filter_inst_lpf_q_pair1_27_8_port, 
      lpf_filter_inst_lpf_q_pair1_27_9_port, 
      lpf_filter_inst_lpf_q_pair1_27_10_port, 
      lpf_filter_inst_lpf_q_pair1_27_11_port, 
      lpf_filter_inst_lpf_q_pair1_27_12_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_0_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_1_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_2_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_3_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_4_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_5_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_6_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_7_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_8_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_9_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_10_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_11_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_12_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_13_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_14_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_15_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_16_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_17_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_18_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_19_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_20_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_21_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_22_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_23_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_24_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_25_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_26_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_27_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_28_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_29_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_30_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_31_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_32_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_33_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_34_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_35_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_36_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_37_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_38_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_39_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_40_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_41_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_42_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_43_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_44_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_45_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_46_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_47_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_48_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_49_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_50_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_51_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_52_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_53_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_54_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_55_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_56_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_57_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_58_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_59_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_60_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_61_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_62_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_63_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_64_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_65_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_66_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_67_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_68_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_69_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_70_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_71_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_72_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_73_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_74_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_75_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_76_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_77_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_78_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_79_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_80_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_81_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_82_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_83_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_84_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_85_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_86_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_87_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_88_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_89_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_90_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_91_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_92_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_93_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_94_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_95_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_96_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_97_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_98_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_99_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_100_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_101_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_102_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_103_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_104_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_105_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_106_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_107_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_108_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_109_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_110_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_111_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_112_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_113_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_114_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_115_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_116_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_117_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_118_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_119_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_120_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_121_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_122_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_123_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_124_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_125_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_126_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_127_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_128_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_129_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_130_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_131_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_132_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_133_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_134_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_135_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_136_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_137_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_138_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_139_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_140_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_141_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_142_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_143_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_144_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_145_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_146_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_147_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_148_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_149_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_150_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_151_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_152_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_153_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_154_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_155_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_156_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_157_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_158_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_159_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_160_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_161_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_162_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_163_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_164_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_165_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_166_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_167_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_168_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_169_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_170_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_171_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_172_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_173_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_174_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_175_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_176_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_177_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_178_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_179_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_180_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_181_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_182_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_183_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_184_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_185_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_186_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_187_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_188_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_189_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_190_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_191_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_192_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_193_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_194_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_195_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_196_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_197_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_198_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_199_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_200_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_201_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_202_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_203_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_204_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_205_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_206_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_207_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_208_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_209_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_210_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_211_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_212_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_213_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_214_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_215_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_216_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_217_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_218_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_219_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_220_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_221_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_222_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_223_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_224_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_225_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_226_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_227_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_228_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_229_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_230_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_231_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_232_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_233_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_234_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_235_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_236_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_237_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_238_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_239_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_240_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_241_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_242_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_243_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_244_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_245_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_246_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_247_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_248_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_249_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_250_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_251_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_252_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_253_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_254_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_255_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_256_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_257_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_258_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_259_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_260_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_261_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_262_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_263_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_264_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_265_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_266_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_267_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_268_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_269_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_270_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_271_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_272_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_273_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_274_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_275_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_276_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_277_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_278_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_279_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_280_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_281_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_282_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_283_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_284_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_285_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_286_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_287_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_288_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_289_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_290_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_291_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_292_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_293_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_294_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_295_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_296_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_297_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_298_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_299_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_300_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_301_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_302_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_303_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_304_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_305_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_306_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_307_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_308_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_309_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_310_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_311_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_312_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_313_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_314_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_315_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_316_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_317_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_318_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_319_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_320_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_321_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_322_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_323_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_324_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_325_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_326_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_327_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_328_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_329_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_330_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_331_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_332_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_333_port, 
      lpf_filter_inst_lpf_q_arx_input_reg_334_port, 
      lpf_filter_inst_lpf_q_add_273_n_1321, lpf_filter_inst_lpf_q_add_273_n1, 
      lpf_filter_inst_lpf_q_add_273_carry_2_port, 
      lpf_filter_inst_lpf_q_add_273_carry_3_port, 
      lpf_filter_inst_lpf_q_add_273_carry_4_port, 
      lpf_filter_inst_lpf_q_add_273_carry_5_port, 
      lpf_filter_inst_lpf_q_add_273_carry_6_port, 
      lpf_filter_inst_lpf_q_add_273_carry_7_port, 
      lpf_filter_inst_lpf_q_add_273_carry_8_port, 
      lpf_filter_inst_lpf_q_add_273_carry_9_port, 
      lpf_filter_inst_lpf_q_add_273_carry_10_port, 
      lpf_filter_inst_lpf_q_add_273_carry_11_port, 
      lpf_filter_inst_lpf_q_add_273_carry_12_port, 
      lpf_filter_inst_lpf_q_add_272_n1, 
      lpf_filter_inst_lpf_q_add_272_carry_2_port, 
      lpf_filter_inst_lpf_q_add_272_carry_3_port, 
      lpf_filter_inst_lpf_q_add_272_carry_4_port, 
      lpf_filter_inst_lpf_q_add_272_carry_5_port, 
      lpf_filter_inst_lpf_q_add_272_carry_6_port, 
      lpf_filter_inst_lpf_q_add_272_carry_7_port, 
      lpf_filter_inst_lpf_q_add_272_carry_8_port, 
      lpf_filter_inst_lpf_q_add_272_carry_9_port, 
      lpf_filter_inst_lpf_q_add_272_carry_10_port, 
      lpf_filter_inst_lpf_q_add_272_carry_11_port, 
      lpf_filter_inst_lpf_q_add_272_carry_12_port, 
      lpf_filter_inst_lpf_q_add_271_n_1316, lpf_filter_inst_lpf_q_add_271_n1, 
      lpf_filter_inst_lpf_q_add_271_carry_2_port, 
      lpf_filter_inst_lpf_q_add_271_carry_3_port, 
      lpf_filter_inst_lpf_q_add_271_carry_4_port, 
      lpf_filter_inst_lpf_q_add_271_carry_5_port, 
      lpf_filter_inst_lpf_q_add_271_carry_6_port, 
      lpf_filter_inst_lpf_q_add_271_carry_7_port, 
      lpf_filter_inst_lpf_q_add_271_carry_8_port, 
      lpf_filter_inst_lpf_q_add_271_carry_9_port, 
      lpf_filter_inst_lpf_q_add_271_carry_10_port, 
      lpf_filter_inst_lpf_q_add_271_carry_11_port, 
      lpf_filter_inst_lpf_q_add_271_carry_12_port, 
      lpf_filter_inst_lpf_q_add_268_n1, 
      lpf_filter_inst_lpf_q_add_268_carry_2_port, 
      lpf_filter_inst_lpf_q_add_268_carry_3_port, 
      lpf_filter_inst_lpf_q_add_268_carry_4_port, 
      lpf_filter_inst_lpf_q_add_268_carry_5_port, 
      lpf_filter_inst_lpf_q_add_268_carry_6_port, 
      lpf_filter_inst_lpf_q_add_268_carry_7_port, 
      lpf_filter_inst_lpf_q_add_268_carry_8_port, 
      lpf_filter_inst_lpf_q_add_268_carry_9_port, 
      lpf_filter_inst_lpf_q_add_268_carry_10_port, 
      lpf_filter_inst_lpf_q_add_268_carry_11_port, 
      lpf_filter_inst_lpf_q_add_268_carry_12_port, 
      lpf_filter_inst_lpf_q_add_264_n_1311, lpf_filter_inst_lpf_q_add_264_n1, 
      lpf_filter_inst_lpf_q_add_264_carry_2_port, 
      lpf_filter_inst_lpf_q_add_264_carry_3_port, 
      lpf_filter_inst_lpf_q_add_264_carry_4_port, 
      lpf_filter_inst_lpf_q_add_264_carry_5_port, 
      lpf_filter_inst_lpf_q_add_264_carry_6_port, 
      lpf_filter_inst_lpf_q_add_264_carry_7_port, 
      lpf_filter_inst_lpf_q_add_264_carry_8_port, 
      lpf_filter_inst_lpf_q_add_264_carry_9_port, 
      lpf_filter_inst_lpf_q_add_264_carry_10_port, 
      lpf_filter_inst_lpf_q_add_264_carry_11_port, 
      lpf_filter_inst_lpf_q_add_264_carry_12_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_n1, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_2_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_q_add_5_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_n1, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_q_add_4_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_n_1079, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_n1, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_q_add_7_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_n_1089, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_n1, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_q_add_8_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_n_1098, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_n1, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_q_add_6_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_n_1104, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_n1, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_23_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n_1109, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n16, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n15, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n14, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n13, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n12, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n11, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n10, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n9, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n8, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n7, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n6, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n5, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n4, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n3, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n1, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_23_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_n_1113, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_n1, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_3_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_4_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_5_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_6_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_7_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_8_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_9_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_10_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_11_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_23_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n_1128, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n29, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n28, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n27, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n26, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n25, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n24, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n23, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n22, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n21, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n20, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n19, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n18, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n17, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n16, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n15, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n14, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n13, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n12, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n11, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n10, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n9, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n8, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n7, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n6, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n5, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n4, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n3, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n2, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_12_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_13_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_14_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_15_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_16_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_17_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_18_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_19_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_20_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_21_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_22_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_23_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_n_1158, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_n1, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_8_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_9_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_10_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_11_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_12_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_13_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_14_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_15_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_16_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_17_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_18_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_285_carry_19_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_n_1268, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_n1, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_2_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_3_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_4_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_5_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_6_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_7_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_8_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_9_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_10_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_11_port, 
      lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_12_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_n_1271, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_n1, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_2_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_3_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_4_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_5_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_6_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_7_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_8_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_9_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_10_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_11_port, 
      lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_12_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_n_1274, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_n1, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_2_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_3_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_4_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_5_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_6_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_7_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_8_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_9_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_10_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_11_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_12_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_13_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n_1279, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n15, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n14, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n13, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n12, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n11, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n10, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n9, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n8, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n7, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n6, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n5, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n4, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n3, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n2, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_n1, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_3_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_4_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_5_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_6_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_7_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_8_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_9_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_10_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_11_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_12_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_13_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_14_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_15_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_16_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_n_1208, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_n1, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_7_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_8_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_9_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_10_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_11_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_12_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_13_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_14_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_15_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_16_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_286_carry_17_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n_1214, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n20, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n19, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n18, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n17, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n16, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n15, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n14, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n13, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n12, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n11, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n10, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n9, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n8, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n7, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n6, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n5, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n4, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n3, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n2, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_n1, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_4_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_5_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_6_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_7_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_8_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_9_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_10_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_11_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_12_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_13_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_14_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_15_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_16_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_17_port, 
      lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_18_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_n_1290, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_n1, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_2_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_3_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_4_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_5_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_6_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_7_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_8_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_9_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_10_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_11_port, 
      lpf_filter_inst_lpf_q_add_1_root_add_277_carry_12_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_n_1293, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_n1, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_2_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_3_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_4_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_5_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_6_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_7_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_8_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_9_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_10_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_11_port, 
      lpf_filter_inst_lpf_q_add_2_root_add_277_carry_12_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_n1, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_2_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_3_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_4_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_5_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_6_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_7_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_8_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_9_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_10_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_11_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_12_port, 
      lpf_filter_inst_lpf_q_add_0_root_add_277_carry_13_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_n_1189, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_n1, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_2_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_3_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_4_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_5_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_6_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_7_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_8_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_9_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_10_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_11_port, 
      lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_12_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n_1194, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n14, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n13, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n12, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n11, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n10, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n9, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n8, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n7, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n6, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n5, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n4, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n3, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n2, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_n1, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_3_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_4_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_5_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_6_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_7_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_8_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_9_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_10_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_11_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_12_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_13_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_14_port, 
      lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_15_port, 
      dam_demodulator_inst_n_1427, dam_demodulator_inst_n_1426, 
      dam_demodulator_inst_n_1425, dam_demodulator_inst_n10, 
      dam_demodulator_inst_n9, dam_demodulator_inst_n8, dam_demodulator_inst_n7
      , dam_demodulator_inst_n6, dam_demodulator_inst_n5, 
      dam_demodulator_inst_n1, dam_demodulator_inst_prod_i_qd_0, 
      dam_demodulator_inst_prod_i_qd_1, dam_demodulator_inst_prod_i_qd_2, 
      dam_demodulator_inst_prod_i_qd_3, dam_demodulator_inst_prod_i_qd_4, 
      dam_demodulator_inst_prod_i_qd_5, dam_demodulator_inst_prod_i_qd_6, 
      dam_demodulator_inst_prod_i_qd_7, dam_demodulator_inst_prod_i_qd_8, 
      dam_demodulator_inst_prod_i_qd_9, dam_demodulator_inst_prod_q_id_0, 
      dam_demodulator_inst_prod_q_id_1, dam_demodulator_inst_prod_q_id_2, 
      dam_demodulator_inst_prod_q_id_3, dam_demodulator_inst_prod_q_id_4, 
      dam_demodulator_inst_prod_q_id_5, dam_demodulator_inst_prod_q_id_6, 
      dam_demodulator_inst_prod_q_id_7, dam_demodulator_inst_prod_q_id_8, 
      dam_demodulator_inst_prod_q_id_9, dam_demodulator_inst_n4, 
      dam_demodulator_inst_n3, dam_demodulator_inst_n2, 
      dam_demodulator_inst_result_2_port, dam_demodulator_inst_result_3_port, 
      dam_demodulator_inst_result_4_port, dam_demodulator_inst_result_5_port, 
      dam_demodulator_inst_result_6_port, dam_demodulator_inst_result_7_port, 
      dam_demodulator_inst_result_8_port, dam_demodulator_inst_result_9_port, 
      dam_demodulator_inst_result_10_port, 
      dam_demodulator_inst_arx_result_reg_2_port, 
      dam_demodulator_inst_arx_result_reg_3_port, 
      dam_demodulator_inst_arx_result_reg_4_port, 
      dam_demodulator_inst_arx_result_reg_5_port, 
      dam_demodulator_inst_arx_result_reg_6_port, 
      dam_demodulator_inst_arx_result_reg_7_port, 
      dam_demodulator_inst_arx_result_reg_8_port, 
      dam_demodulator_inst_arx_result_reg_9_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_0_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_1_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_2_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_3_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_4_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_5_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_6_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_7_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_8_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_9_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_10_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_11_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_12_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_13_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_14_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_15_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_16_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_17_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_18_port, 
      dam_demodulator_inst_arx_dem_samples_q_reg_19_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_0_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_1_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_2_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_3_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_4_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_5_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_6_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_7_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_8_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_9_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_10_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_11_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_12_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_13_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_14_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_15_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_16_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_17_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_18_port, 
      dam_demodulator_inst_arx_dem_samples_i_reg_19_port, 
      dam_demodulator_inst_mult_131_n101, dam_demodulator_inst_mult_131_n100, 
      dam_demodulator_inst_mult_131_n99, dam_demodulator_inst_mult_131_n98, 
      dam_demodulator_inst_mult_131_n97, dam_demodulator_inst_mult_131_n96, 
      dam_demodulator_inst_mult_131_n95, dam_demodulator_inst_mult_131_n94, 
      dam_demodulator_inst_mult_131_n93, dam_demodulator_inst_mult_131_n92, 
      dam_demodulator_inst_mult_131_n56, dam_demodulator_inst_mult_131_n55, 
      dam_demodulator_inst_mult_131_n54, dam_demodulator_inst_mult_131_n53, 
      dam_demodulator_inst_mult_131_n52, dam_demodulator_inst_mult_131_n51, 
      dam_demodulator_inst_mult_131_n50, dam_demodulator_inst_mult_131_n49, 
      dam_demodulator_inst_mult_131_n48, dam_demodulator_inst_mult_131_n47, 
      dam_demodulator_inst_mult_131_n46, dam_demodulator_inst_mult_131_n45, 
      dam_demodulator_inst_mult_131_n43, dam_demodulator_inst_mult_131_n42, 
      dam_demodulator_inst_mult_131_n41, dam_demodulator_inst_mult_131_n39, 
      dam_demodulator_inst_mult_131_n38, dam_demodulator_inst_mult_131_n37, 
      dam_demodulator_inst_mult_131_n36, dam_demodulator_inst_mult_131_n35, 
      dam_demodulator_inst_mult_131_n34, dam_demodulator_inst_mult_131_n33, 
      dam_demodulator_inst_mult_131_n32, dam_demodulator_inst_mult_131_n31, 
      dam_demodulator_inst_mult_131_n30, dam_demodulator_inst_mult_131_n29, 
      dam_demodulator_inst_mult_131_n28, dam_demodulator_inst_mult_131_n27, 
      dam_demodulator_inst_mult_131_n26, dam_demodulator_inst_mult_131_n25, 
      dam_demodulator_inst_mult_131_n24, dam_demodulator_inst_mult_131_n23, 
      dam_demodulator_inst_mult_131_n22, dam_demodulator_inst_mult_131_n21, 
      dam_demodulator_inst_mult_131_n20, dam_demodulator_inst_mult_131_n19, 
      dam_demodulator_inst_mult_131_n18, dam_demodulator_inst_mult_131_n17, 
      dam_demodulator_inst_mult_131_n16, dam_demodulator_inst_mult_131_n15, 
      dam_demodulator_inst_mult_131_n14, dam_demodulator_inst_mult_131_n13, 
      dam_demodulator_inst_mult_131_n12, dam_demodulator_inst_mult_131_n11, 
      dam_demodulator_inst_mult_131_n10, dam_demodulator_inst_mult_131_n9, 
      dam_demodulator_inst_mult_131_n8, dam_demodulator_inst_mult_131_n7, 
      dam_demodulator_inst_mult_131_n6, dam_demodulator_inst_mult_131_n5, 
      dam_demodulator_inst_mult_131_n4, dam_demodulator_inst_mult_131_n3, 
      dam_demodulator_inst_mult_131_n2, dam_demodulator_inst_mult_131_n1, 
      dam_demodulator_inst_mult_130_n101, dam_demodulator_inst_mult_130_n100, 
      dam_demodulator_inst_mult_130_n99, dam_demodulator_inst_mult_130_n98, 
      dam_demodulator_inst_mult_130_n97, dam_demodulator_inst_mult_130_n96, 
      dam_demodulator_inst_mult_130_n95, dam_demodulator_inst_mult_130_n94, 
      dam_demodulator_inst_mult_130_n93, dam_demodulator_inst_mult_130_n92, 
      dam_demodulator_inst_mult_130_n56, dam_demodulator_inst_mult_130_n55, 
      dam_demodulator_inst_mult_130_n54, dam_demodulator_inst_mult_130_n53, 
      dam_demodulator_inst_mult_130_n52, dam_demodulator_inst_mult_130_n51, 
      dam_demodulator_inst_mult_130_n50, dam_demodulator_inst_mult_130_n49, 
      dam_demodulator_inst_mult_130_n48, dam_demodulator_inst_mult_130_n47, 
      dam_demodulator_inst_mult_130_n46, dam_demodulator_inst_mult_130_n45, 
      dam_demodulator_inst_mult_130_n43, dam_demodulator_inst_mult_130_n42, 
      dam_demodulator_inst_mult_130_n41, dam_demodulator_inst_mult_130_n39, 
      dam_demodulator_inst_mult_130_n38, dam_demodulator_inst_mult_130_n37, 
      dam_demodulator_inst_mult_130_n36, dam_demodulator_inst_mult_130_n35, 
      dam_demodulator_inst_mult_130_n34, dam_demodulator_inst_mult_130_n33, 
      dam_demodulator_inst_mult_130_n32, dam_demodulator_inst_mult_130_n31, 
      dam_demodulator_inst_mult_130_n30, dam_demodulator_inst_mult_130_n29, 
      dam_demodulator_inst_mult_130_n28, dam_demodulator_inst_mult_130_n27, 
      dam_demodulator_inst_mult_130_n26, dam_demodulator_inst_mult_130_n25, 
      dam_demodulator_inst_mult_130_n24, dam_demodulator_inst_mult_130_n23, 
      dam_demodulator_inst_mult_130_n22, dam_demodulator_inst_mult_130_n21, 
      dam_demodulator_inst_mult_130_n20, dam_demodulator_inst_mult_130_n19, 
      dam_demodulator_inst_mult_130_n18, dam_demodulator_inst_mult_130_n17, 
      dam_demodulator_inst_mult_130_n16, dam_demodulator_inst_mult_130_n15, 
      dam_demodulator_inst_mult_130_n14, dam_demodulator_inst_mult_130_n13, 
      dam_demodulator_inst_mult_130_n12, dam_demodulator_inst_mult_130_n11, 
      dam_demodulator_inst_mult_130_n10, dam_demodulator_inst_mult_130_n9, 
      dam_demodulator_inst_mult_130_n8, dam_demodulator_inst_mult_130_n7, 
      dam_demodulator_inst_mult_130_n6, dam_demodulator_inst_mult_130_n5, 
      dam_demodulator_inst_mult_130_n4, dam_demodulator_inst_mult_130_n3, 
      dam_demodulator_inst_mult_130_n2, dam_demodulator_inst_mult_130_n1, 
      dam_demodulator_inst_sub_132_n_1004, dam_demodulator_inst_sub_132_n11, 
      dam_demodulator_inst_sub_132_n10, dam_demodulator_inst_sub_132_n9, 
      dam_demodulator_inst_sub_132_n8, dam_demodulator_inst_sub_132_n7, 
      dam_demodulator_inst_sub_132_n6, dam_demodulator_inst_sub_132_n5, 
      dam_demodulator_inst_sub_132_n4, dam_demodulator_inst_sub_132_n3, 
      dam_demodulator_inst_sub_132_n2, dam_demodulator_inst_sub_132_n1, 
      dam_demodulator_inst_sub_132_carry_2_port, 
      dam_demodulator_inst_sub_132_carry_3_port, 
      dam_demodulator_inst_sub_132_carry_4_port, 
      dam_demodulator_inst_sub_132_carry_5_port, 
      dam_demodulator_inst_sub_132_carry_6_port, 
      dam_demodulator_inst_sub_132_carry_7_port, 
      dam_demodulator_inst_sub_132_carry_8_port, 
      dam_demodulator_inst_sub_132_carry_9_port, 
      dam_demodulator_inst_sub_132_carry_10_port, sl_slicer_inst_n_1424, 
      sl_slicer_inst_n_1423, sl_slicer_inst_n_1422, sl_slicer_inst_n101, 
      sl_slicer_inst_n9, sl_slicer_inst_n8, sl_slicer_inst_n7, 
      sl_slicer_inst_n6, sl_slicer_inst_n100, sl_slicer_inst_sum0_1_0, 
      sl_slicer_inst_sum0_1_1, sl_slicer_inst_sum0_1_2, sl_slicer_inst_sum0_1_3
      , sl_slicer_inst_sum0_1_4, sl_slicer_inst_sum0_1_5, 
      sl_slicer_inst_sum0_1_6, sl_slicer_inst_sum0_1_7, sl_slicer_inst_sum2_3_0
      , sl_slicer_inst_sum2_3_1, sl_slicer_inst_sum2_3_2, 
      sl_slicer_inst_sum2_3_3, sl_slicer_inst_sum2_3_4, sl_slicer_inst_sum2_3_5
      , sl_slicer_inst_sum2_3_6, sl_slicer_inst_sum2_3_7, sl_slicer_inst_n5, 
      sl_slicer_inst_n4, sl_slicer_inst_n3, sl_slicer_inst_n2, 
      sl_slicer_inst_N1, sl_slicer_inst_counter_1, 
      sl_slicer_inst_sum0_1_2_3_0_port, sl_slicer_inst_sum0_1_2_3_1_port, 
      sl_slicer_inst_sum0_1_2_3_2_port, sl_slicer_inst_sum0_1_2_3_3_port, 
      sl_slicer_inst_sum0_1_2_3_4_port, sl_slicer_inst_sum0_1_2_3_5_port, 
      sl_slicer_inst_sum0_1_2_3_6_port, sl_slicer_inst_sum0_1_2_3_7_port, 
      sl_slicer_inst_sum0_1_2_3_8_port, sl_slicer_inst_arx_counter_reg_0_port, 
      sl_slicer_inst_arx_counter_reg_1_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_0_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_1_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_2_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_3_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_4_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_5_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_6_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_7_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_8_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_9_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_10_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_11_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_12_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_13_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_14_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_15_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_16_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_17_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_18_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_19_port, 
      sl_slicer_inst_arx_slicer_fifo_reg_20_port, 
      sl_slicer_inst_add_2_root_add_122_n_1217, 
      sl_slicer_inst_add_2_root_add_122_n1, 
      sl_slicer_inst_add_2_root_add_122_carry_2_port, 
      sl_slicer_inst_add_2_root_add_122_carry_3_port, 
      sl_slicer_inst_add_2_root_add_122_carry_4_port, 
      sl_slicer_inst_add_2_root_add_122_carry_5_port, 
      sl_slicer_inst_add_2_root_add_122_carry_6_port, 
      sl_slicer_inst_add_2_root_add_122_carry_7_port, 
      sl_slicer_inst_add_1_root_add_122_n_1220, 
      sl_slicer_inst_add_1_root_add_122_n1, 
      sl_slicer_inst_add_1_root_add_122_carry_2_port, 
      sl_slicer_inst_add_1_root_add_122_carry_3_port, 
      sl_slicer_inst_add_1_root_add_122_carry_4_port, 
      sl_slicer_inst_add_1_root_add_122_carry_5_port, 
      sl_slicer_inst_add_1_root_add_122_carry_6_port, 
      sl_slicer_inst_add_1_root_add_122_carry_7_port, 
      sl_slicer_inst_add_0_root_add_122_n_1223, 
      sl_slicer_inst_add_0_root_add_122_n1, 
      sl_slicer_inst_add_0_root_add_122_carry_2_port, 
      sl_slicer_inst_add_0_root_add_122_carry_3_port, 
      sl_slicer_inst_add_0_root_add_122_carry_4_port, 
      sl_slicer_inst_add_0_root_add_122_carry_5_port, 
      sl_slicer_inst_add_0_root_add_122_carry_6_port, 
      sl_slicer_inst_add_0_root_add_122_carry_7_port, 
      sl_slicer_inst_add_0_root_add_122_carry_8_port : std_logic;

begin
   slicer_out <= slicer_out_port;
   
   U3 : TIEHI port map( Z => n_Logic1);
   U4 : TIELO port map( Z => n_Logic0);
   cg_U4 : AND2D1 port map( A1 => cg_counter_1_port, A2 => cg_counter_0_port, Z
                           => cg_N2);
   cg_U3 : INVD1 port map( A => cg_counter_0_port, Z => cg_n10);
   cg_counter_reg_0 : DFFRPQ1 port map( D => cg_n10, CK => clk, RB => rstn, Q 
                           => cg_counter_0_port);
   cg_counter_reg_1 : DFFRPQ1 port map( D => cg_N1, CK => clk, RB => rstn, Q =>
                           cg_counter_1_port);
   cg_clk4_reg : DFFRPQ1 port map( D => cg_N2, CK => clk, RB => rstn, Q => clk4
                           );
   cg_U5 : EXNOR2D1 port map( A1 => cg_counter_1_port, A2 => cg_n10, Z => cg_N1
                           );
   mx_mixer_inst_U136 : EXOR2D1 port map( A1 => mx_mixer_inst_n77, A2 => 
                           mx_mixer_inst_n76, Z => mx_mixer_inst_N58);
   mx_mixer_inst_U135 : AND2D1 port map( A1 => mx_mixer_inst_n76, A2 => 
                           mx_mixer_inst_n77, Z => 
                           mx_mixer_inst_r377_carry_8_port);
   mx_mixer_inst_U134 : EXOR2D1 port map( A1 => mx_mixer_inst_n78, A2 => 
                           mx_mixer_inst_r377_carry_8_port, Z => 
                           mx_mixer_inst_N59);
   mx_mixer_inst_U133 : AND2D1 port map( A1 => mx_mixer_inst_r377_carry_8_port,
                           A2 => mx_mixer_inst_n78, Z => 
                           mx_mixer_inst_r377_carry_9_port);
   mx_mixer_inst_U132 : EXOR2D1 port map( A1 => mx_mixer_inst_n79, A2 => 
                           mx_mixer_inst_r377_carry_9_port, Z => 
                           mx_mixer_inst_N60);
   mx_mixer_inst_U131 : AND2D1 port map( A1 => mx_mixer_inst_r377_carry_9_port,
                           A2 => mx_mixer_inst_n79, Z => 
                           mx_mixer_inst_r377_carry_10_port);
   mx_mixer_inst_U130 : EXOR2D1 port map( A1 => mx_mixer_inst_n80, A2 => 
                           mx_mixer_inst_r377_carry_10_port, Z => 
                           mx_mixer_inst_N61);
   mx_mixer_inst_U129 : AND2D1 port map( A1 => mx_mixer_inst_r377_carry_10_port
                           , A2 => mx_mixer_inst_n80, Z => 
                           mx_mixer_inst_r377_carry_11_port);
   mx_mixer_inst_U128 : EXOR2D1 port map( A1 => mx_mixer_inst_n81, A2 => 
                           mx_mixer_inst_r377_carry_11_port, Z => 
                           mx_mixer_inst_N62);
   mx_mixer_inst_U127 : AND2D1 port map( A1 => mx_mixer_inst_r377_carry_11_port
                           , A2 => mx_mixer_inst_n81, Z => 
                           mx_mixer_inst_r377_carry_12_port);
   mx_mixer_inst_U126 : EXOR2D1 port map( A1 => mx_mixer_inst_n82, A2 => 
                           mx_mixer_inst_r377_carry_12_port, Z => 
                           mx_mixer_inst_N63);
   mx_mixer_inst_U125 : AND2D1 port map( A1 => mx_mixer_inst_r377_carry_12_port
                           , A2 => mx_mixer_inst_n82, Z => 
                           mx_mixer_inst_r377_carry_13_port);
   mx_mixer_inst_U124 : EXOR2D1 port map( A1 => mx_mixer_inst_n83, A2 => 
                           mx_mixer_inst_r377_carry_13_port, Z => 
                           mx_mixer_inst_N64);
   mx_mixer_inst_U123 : AND2D1 port map( A1 => mx_mixer_inst_r377_carry_13_port
                           , A2 => mx_mixer_inst_n83, Z => 
                           mx_mixer_inst_r377_carry_14_port);
   mx_mixer_inst_U122 : EXOR2D1 port map( A1 => mx_mixer_inst_n84, A2 => 
                           mx_mixer_inst_r377_carry_14_port, Z => 
                           mx_mixer_inst_N65);
   mx_mixer_inst_U121 : AND2D1 port map( A1 => mx_mixer_inst_r377_carry_14_port
                           , A2 => mx_mixer_inst_n84, Z => 
                           mx_mixer_inst_r377_carry_15_port);
   mx_mixer_inst_U120 : EXOR2D1 port map( A1 => mx_mixer_inst_n85, A2 => 
                           mx_mixer_inst_r377_carry_15_port, Z => 
                           mx_mixer_inst_N66);
   mx_mixer_inst_U119 : AND2D1 port map( A1 => mx_mixer_inst_r377_carry_15_port
                           , A2 => mx_mixer_inst_n85, Z => 
                           mx_mixer_inst_r377_carry_16_port);
   mx_mixer_inst_U118 : EXOR2D1 port map( A1 => mx_mixer_inst_n86, A2 => 
                           mx_mixer_inst_r377_carry_16_port, Z => 
                           mx_mixer_inst_N67);
   mx_mixer_inst_U117 : NAN2D1 port map( A1 => mx_mixer_inst_n610, A2 => 
                           mx_mixer_inst_n600, Z => mixer_out_q_11_port);
   mx_mixer_inst_U116 : AOI22D1 port map( A1 => mx_mixer_inst_N68, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N44, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n600);
   mx_mixer_inst_U115 : AOI22D1 port map( A1 => mixer_in(11), A2 => 
                           mx_mixer_inst_n570, B1 => mixer_in(11), B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n610);
   mx_mixer_inst_U114 : NAN2D1 port map( A1 => mx_mixer_inst_n550, A2 => 
                           mx_mixer_inst_n540, Z => mixer_out_q_10_port);
   mx_mixer_inst_U113 : AOI22D1 port map( A1 => mx_mixer_inst_N67, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N43, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n540);
   mx_mixer_inst_U112 : AOI22D1 port map( A1 => mixer_in(10), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N55, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n550);
   mx_mixer_inst_U111 : NAN2D1 port map( A1 => mx_mixer_inst_n530, A2 => 
                           mx_mixer_inst_n520, Z => mixer_out_q_9_port);
   mx_mixer_inst_U110 : AOI22D1 port map( A1 => mx_mixer_inst_N66, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N42, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n520);
   mx_mixer_inst_U109 : AOI22D1 port map( A1 => mixer_in(9), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N54, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n530);
   mx_mixer_inst_U108 : NAN2D1 port map( A1 => mx_mixer_inst_n510, A2 => 
                           mx_mixer_inst_n500, Z => mixer_out_q_8_port);
   mx_mixer_inst_U107 : AOI22D1 port map( A1 => mx_mixer_inst_N65, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N41, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n500);
   mx_mixer_inst_U106 : AOI22D1 port map( A1 => mixer_in(8), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N53, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n510);
   mx_mixer_inst_U105 : NAN2D1 port map( A1 => mx_mixer_inst_n490, A2 => 
                           mx_mixer_inst_n480, Z => mixer_out_q_7_port);
   mx_mixer_inst_U104 : AOI22D1 port map( A1 => mx_mixer_inst_N64, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N40, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n480);
   mx_mixer_inst_U103 : AOI22D1 port map( A1 => mixer_in(7), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N52, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n490);
   mx_mixer_inst_U102 : NAN2D1 port map( A1 => mx_mixer_inst_n470, A2 => 
                           mx_mixer_inst_n460, Z => mixer_out_q_6_port);
   mx_mixer_inst_U101 : AOI22D1 port map( A1 => mx_mixer_inst_N63, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N39, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n460);
   mx_mixer_inst_U100 : AOI22D1 port map( A1 => mixer_in(6), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N51, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n470);
   mx_mixer_inst_U99 : NAN2D1 port map( A1 => mx_mixer_inst_n450, A2 => 
                           mx_mixer_inst_n440, Z => mixer_out_q_5_port);
   mx_mixer_inst_U98 : AOI22D1 port map( A1 => mx_mixer_inst_N62, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N38, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n440);
   mx_mixer_inst_U97 : AOI22D1 port map( A1 => mixer_in(5), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N50, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n450);
   mx_mixer_inst_U96 : NAN2D1 port map( A1 => mx_mixer_inst_n430, A2 => 
                           mx_mixer_inst_n420, Z => mixer_out_q_4_port);
   mx_mixer_inst_U95 : AOI22D1 port map( A1 => mx_mixer_inst_N61, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N37, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n420);
   mx_mixer_inst_U94 : AOI22D1 port map( A1 => mixer_in(4), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N49, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n430);
   mx_mixer_inst_U93 : NAN2D1 port map( A1 => mx_mixer_inst_n410, A2 => 
                           mx_mixer_inst_n400, Z => mixer_out_q_3_port);
   mx_mixer_inst_U92 : AOI22D1 port map( A1 => mx_mixer_inst_N60, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N36, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n400);
   mx_mixer_inst_U91 : AOI22D1 port map( A1 => mixer_in(3), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N48, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n410);
   mx_mixer_inst_U90 : NAN2D1 port map( A1 => mx_mixer_inst_n390, A2 => 
                           mx_mixer_inst_n380, Z => mixer_out_q_2_port);
   mx_mixer_inst_U89 : AOI22D1 port map( A1 => mx_mixer_inst_N59, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N35, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n380);
   mx_mixer_inst_U88 : AOI22D1 port map( A1 => mixer_in(2), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N47, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n390);
   mx_mixer_inst_U87 : NAN2D1 port map( A1 => mx_mixer_inst_n370, A2 => 
                           mx_mixer_inst_n360, Z => mixer_out_q_1_port);
   mx_mixer_inst_U86 : AOI22D1 port map( A1 => mx_mixer_inst_N58, A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N34, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n360);
   mx_mixer_inst_U85 : AOI22D1 port map( A1 => mixer_in(1), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N46, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n370);
   mx_mixer_inst_U84 : NAN2D1 port map( A1 => mx_mixer_inst_n350, A2 => 
                           mx_mixer_inst_n340, Z => mixer_out_q_0_port);
   mx_mixer_inst_U83 : AOI22D1 port map( A1 => mixer_in(0), A2 => 
                           mx_mixer_inst_n590, B1 => mx_mixer_inst_N33, B2 => 
                           mx_mixer_inst_n580, Z => mx_mixer_inst_n340);
   mx_mixer_inst_U82 : AOI22D1 port map( A1 => mixer_in(0), A2 => 
                           mx_mixer_inst_n570, B1 => mx_mixer_inst_N45, B2 => 
                           mx_mixer_inst_n560, Z => mx_mixer_inst_n350);
   mx_mixer_inst_U81 : AND2D1 port map( A1 => mx_mixer_inst_arx_i_reg_1_port, 
                           A2 => mx_mixer_inst_n75, Z => mx_mixer_inst_n330);
   mx_mixer_inst_U80 : OAI211D1 port map( A1 => mx_mixer_inst_n73, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n31, C => 
                           mx_mixer_inst_n30, Z => mixer_out_i_11_port);
   mx_mixer_inst_U79 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(11), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N68, Z => mx_mixer_inst_n30);
   mx_mixer_inst_U78 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mixer_in(11), Z => mx_mixer_inst_n31);
   mx_mixer_inst_U77 : OAI211D1 port map( A1 => mx_mixer_inst_n72, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n26, C => 
                           mx_mixer_inst_n25, Z => mixer_out_i_10_port);
   mx_mixer_inst_U76 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(10), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N67, Z => mx_mixer_inst_n25);
   mx_mixer_inst_U75 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N55, Z => mx_mixer_inst_n26);
   mx_mixer_inst_U74 : OAI211D1 port map( A1 => mx_mixer_inst_n71, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n24, C => 
                           mx_mixer_inst_n23, Z => mixer_out_i_9_port);
   mx_mixer_inst_U73 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(9), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N66, Z => mx_mixer_inst_n23);
   mx_mixer_inst_U72 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N54, Z => mx_mixer_inst_n24);
   mx_mixer_inst_U71 : OAI211D1 port map( A1 => mx_mixer_inst_n70, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n22, C => 
                           mx_mixer_inst_n21, Z => mixer_out_i_8_port);
   mx_mixer_inst_U70 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(8), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N65, Z => mx_mixer_inst_n21);
   mx_mixer_inst_U69 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N53, Z => mx_mixer_inst_n22);
   mx_mixer_inst_U68 : OAI211D1 port map( A1 => mx_mixer_inst_n69, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n20, C => 
                           mx_mixer_inst_n19, Z => mixer_out_i_7_port);
   mx_mixer_inst_U67 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(7), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N64, Z => mx_mixer_inst_n19);
   mx_mixer_inst_U66 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N52, Z => mx_mixer_inst_n20);
   mx_mixer_inst_U65 : OAI211D1 port map( A1 => mx_mixer_inst_n680, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n18, C => 
                           mx_mixer_inst_n17, Z => mixer_out_i_6_port);
   mx_mixer_inst_U64 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(6), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N63, Z => mx_mixer_inst_n17);
   mx_mixer_inst_U63 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N51, Z => mx_mixer_inst_n18);
   mx_mixer_inst_U62 : OAI211D1 port map( A1 => mx_mixer_inst_n670, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n16, C => 
                           mx_mixer_inst_n15, Z => mixer_out_i_5_port);
   mx_mixer_inst_U61 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(5), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N62, Z => mx_mixer_inst_n15);
   mx_mixer_inst_U60 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N50, Z => mx_mixer_inst_n16);
   mx_mixer_inst_U59 : OAI211D1 port map( A1 => mx_mixer_inst_n660, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n14, C => 
                           mx_mixer_inst_n13, Z => mixer_out_i_4_port);
   mx_mixer_inst_U58 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(4), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N61, Z => mx_mixer_inst_n13);
   mx_mixer_inst_U57 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N49, Z => mx_mixer_inst_n14);
   mx_mixer_inst_U56 : OAI211D1 port map( A1 => mx_mixer_inst_n650, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n12, C => 
                           mx_mixer_inst_n11, Z => mixer_out_i_3_port);
   mx_mixer_inst_U55 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(3), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N60, Z => mx_mixer_inst_n11);
   mx_mixer_inst_U54 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N48, Z => mx_mixer_inst_n12);
   mx_mixer_inst_U53 : OAI211D1 port map( A1 => mx_mixer_inst_n640, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n10, C => 
                           mx_mixer_inst_n9, Z => mixer_out_i_2_port);
   mx_mixer_inst_U52 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(2), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N59, Z => mx_mixer_inst_n9);
   mx_mixer_inst_U51 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N47, Z => mx_mixer_inst_n10);
   mx_mixer_inst_U50 : OAI211D1 port map( A1 => mx_mixer_inst_n630, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n8, C => 
                           mx_mixer_inst_n7, Z => mixer_out_i_1_port);
   mx_mixer_inst_U49 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(1), B1 => mx_mixer_inst_n28, B2 => 
                           mx_mixer_inst_N58, Z => mx_mixer_inst_n7);
   mx_mixer_inst_U48 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N46, Z => mx_mixer_inst_n8);
   mx_mixer_inst_U47 : OAI211D1 port map( A1 => mx_mixer_inst_n620, A2 => 
                           mx_mixer_inst_n32, B => mx_mixer_inst_n6, C => 
                           mx_mixer_inst_n5, Z => mixer_out_i_0_port);
   mx_mixer_inst_U46 : AOI22D1 port map( A1 => mx_mixer_inst_n29, A2 => 
                           mixer_in(0), B1 => mx_mixer_inst_n28, B2 => 
                           mixer_in(0), Z => mx_mixer_inst_n5);
   mx_mixer_inst_U45 : NOR2D1 port map( A1 => mx_mixer_inst_arx_i_reg_0_port, 
                           A2 => mx_mixer_inst_arx_i_reg_1_port, Z => 
                           mx_mixer_inst_n4);
   mx_mixer_inst_U44 : NAN2D1 port map( A1 => mx_mixer_inst_n27, A2 => 
                           mx_mixer_inst_N45, Z => mx_mixer_inst_n6);
   mx_mixer_inst_U43 : EXOR2D1 port map( A1 => mx_mixer_inst_arx_i_reg_1_port, 
                           A2 => mx_mixer_inst_arx_i_reg_2_port, Z => 
                           mx_mixer_inst_n3);
   mx_mixer_inst_U42 : TIEHI port map( Z => mx_mixer_inst_n87);
   mx_mixer_inst_U41 : TIELO port map( Z => mx_mixer_inst_n88);
   mx_mixer_inst_U40 : NAN2D1 port map( A1 => mx_mixer_inst_arx_i_reg_1_port, 
                           A2 => mx_mixer_inst_arx_i_reg_0_port, Z => 
                           mx_mixer_inst_n2);
   mx_mixer_inst_U39 : EXNOR2D1 port map( A1 => mx_mixer_inst_arx_i_reg_2_port,
                           A2 => mx_mixer_inst_n2, Z => mx_mixer_inst_i_2_port)
                           ;
   mx_mixer_inst_U38 : NOR2D1 port map( A1 => mx_mixer_inst_n75, A2 => 
                           mx_mixer_inst_arx_i_reg_2_port, Z => 
                           mx_mixer_inst_n580);
   mx_mixer_inst_U37 : INVD1 port map( A => mx_mixer_inst_arx_i_reg_2_port, Z 
                           => mx_mixer_inst_n74);
   mx_mixer_inst_U36 : NOR2M1D1 port map( A1 => mx_mixer_inst_n4, A2 => 
                           mx_mixer_inst_arx_i_reg_2_port, Z => 
                           mx_mixer_inst_n29);
   mx_mixer_inst_U35 : NAN2D1 port map( A1 => mx_mixer_inst_arx_i_reg_0_port, 
                           A2 => mx_mixer_inst_n3, Z => mx_mixer_inst_n32);
   mx_mixer_inst_U34 : INVD1 port map( A => mx_mixer_inst_arx_i_reg_0_port, Z 
                           => mx_mixer_inst_n75);
   mx_mixer_inst_U33 : NOR2M1D1 port map( A1 => mx_mixer_inst_n330, A2 => 
                           mx_mixer_inst_arx_i_reg_2_port, Z => 
                           mx_mixer_inst_n590);
   mx_mixer_inst_U32 : INVD1 port map( A => mixer_in(10), Z => 
                           mx_mixer_inst_n86);
   mx_mixer_inst_U31 : INVD1 port map( A => mixer_in(9), Z => mx_mixer_inst_n85
                           );
   mx_mixer_inst_U30 : INVD1 port map( A => mixer_in(8), Z => mx_mixer_inst_n84
                           );
   mx_mixer_inst_U29 : INVD1 port map( A => mixer_in(7), Z => mx_mixer_inst_n83
                           );
   mx_mixer_inst_U28 : INVD1 port map( A => mixer_in(6), Z => mx_mixer_inst_n82
                           );
   mx_mixer_inst_U27 : INVD1 port map( A => mixer_in(5), Z => mx_mixer_inst_n81
                           );
   mx_mixer_inst_U26 : INVD1 port map( A => mx_mixer_inst_N33, Z => 
                           mx_mixer_inst_n620);
   mx_mixer_inst_U25 : INVD1 port map( A => mixer_in(4), Z => mx_mixer_inst_n80
                           );
   mx_mixer_inst_U24 : INVD1 port map( A => mx_mixer_inst_N34, Z => 
                           mx_mixer_inst_n630);
   mx_mixer_inst_U23 : INVD1 port map( A => mixer_in(3), Z => mx_mixer_inst_n79
                           );
   mx_mixer_inst_U22 : INVD1 port map( A => mixer_in(2), Z => mx_mixer_inst_n78
                           );
   mx_mixer_inst_U21 : INVD1 port map( A => mx_mixer_inst_N35, Z => 
                           mx_mixer_inst_n640);
   mx_mixer_inst_U20 : INVD1 port map( A => mixer_in(0), Z => mx_mixer_inst_n76
                           );
   mx_mixer_inst_U19 : INVD1 port map( A => mixer_in(1), Z => mx_mixer_inst_n77
                           );
   mx_mixer_inst_U18 : NAN2D1 port map( A1 => mx_mixer_inst_r377_carry_16_port,
                           A2 => mx_mixer_inst_n86, Z => mx_mixer_inst_n1);
   mx_mixer_inst_U17 : EXOR2D1 port map( A1 => mixer_in(11), A2 => 
                           mx_mixer_inst_n1, Z => mx_mixer_inst_N68);
   mx_mixer_inst_U16 : INVD1 port map( A => mx_mixer_inst_N36, Z => 
                           mx_mixer_inst_n650);
   mx_mixer_inst_U15 : INVD1 port map( A => mx_mixer_inst_N37, Z => 
                           mx_mixer_inst_n660);
   mx_mixer_inst_U14 : INVD1 port map( A => mx_mixer_inst_N38, Z => 
                           mx_mixer_inst_n670);
   mx_mixer_inst_U13 : INVD1 port map( A => mx_mixer_inst_N39, Z => 
                           mx_mixer_inst_n680);
   mx_mixer_inst_U12 : INVD1 port map( A => mx_mixer_inst_N40, Z => 
                           mx_mixer_inst_n69);
   mx_mixer_inst_U11 : INVD1 port map( A => mx_mixer_inst_N41, Z => 
                           mx_mixer_inst_n70);
   mx_mixer_inst_U10 : INVD1 port map( A => mx_mixer_inst_N42, Z => 
                           mx_mixer_inst_n71);
   mx_mixer_inst_U9 : INVD1 port map( A => mx_mixer_inst_N43, Z => 
                           mx_mixer_inst_n72);
   mx_mixer_inst_U7 : INVD1 port map( A => mx_mixer_inst_N44, Z => 
                           mx_mixer_inst_n73);
   mx_mixer_inst_U6 : NOR2D1 port map( A1 => mx_mixer_inst_n74, A2 => 
                           mx_mixer_inst_n75, Z => mx_mixer_inst_n560);
   mx_mixer_inst_U5 : NOR2M1D1 port map( A1 => mx_mixer_inst_n4, A2 => 
                           mx_mixer_inst_n74, Z => mx_mixer_inst_n28);
   mx_mixer_inst_U4 : NOR2M1D1 port map( A1 => mx_mixer_inst_n330, A2 => 
                           mx_mixer_inst_n74, Z => mx_mixer_inst_n570);
   mx_mixer_inst_U3 : NOR2D1 port map( A1 => mx_mixer_inst_n3, A2 => 
                           mx_mixer_inst_n75, Z => mx_mixer_inst_n27);
   mx_mixer_inst_arx_i_reg_reg_2 : DFFRPQ1 port map( D => 
                           mx_mixer_inst_i_2_port, CK => clk, RB => rstn, Q => 
                           mx_mixer_inst_arx_i_reg_2_port);
   mx_mixer_inst_arx_i_reg_reg_0 : DFFRPQ1 port map( D => mx_mixer_inst_n75, CK
                           => clk, RB => rstn, Q => 
                           mx_mixer_inst_arx_i_reg_0_port);
   mx_mixer_inst_arx_i_reg_reg_1 : DFFRPQ1 port map( D => 
                           mx_mixer_inst_i_1_port, CK => clk, RB => rstn, Q => 
                           mx_mixer_inst_arx_i_reg_1_port);
   mx_mixer_inst_U8 : EXNOR2D1 port map( A1 => mx_mixer_inst_arx_i_reg_1_port, 
                           A2 => mx_mixer_inst_n75, Z => mx_mixer_inst_i_1_port
                           );
   mx_mixer_inst_r375_U84 : OAI22D1 port map( A1 => mx_mixer_inst_r375_n125, A2
                           => mx_mixer_inst_r375_n124, B1 => 
                           mx_mixer_inst_r375_n125, B2 => 
                           mx_mixer_inst_r375_n126, Z => 
                           mx_mixer_inst_r375_n135);
   mx_mixer_inst_r375_U83 : NAN2D1 port map( A1 => mx_mixer_inst_r375_n135, A2 
                           => mixer_in(3), Z => mx_mixer_inst_r375_n133);
   mx_mixer_inst_r375_U82 : NAN2D1 port map( A1 => mx_mixer_inst_r375_n135, A2 
                           => mixer_in(2), Z => mx_mixer_inst_r375_n134);
   mx_mixer_inst_r375_U81 : OAI211D1 port map( A1 => mx_mixer_inst_r375_n124, 
                           A2 => mx_mixer_inst_r375_n123, B => 
                           mx_mixer_inst_r375_n133, C => 
                           mx_mixer_inst_r375_n134, Z => 
                           mx_mixer_inst_r375_n132);
   mx_mixer_inst_r375_U80 : NAN2D1 port map( A1 => mx_mixer_inst_r375_n53, A2 
                           => mx_mixer_inst_r375_n132, Z => 
                           mx_mixer_inst_r375_n130);
   mx_mixer_inst_r375_U79 : NAN2D1 port map( A1 => mixer_in(0), A2 => 
                           mx_mixer_inst_r375_n132, Z => 
                           mx_mixer_inst_r375_n131);
   mx_mixer_inst_r375_U78 : OAI211D1 port map( A1 => mx_mixer_inst_r375_n126, 
                           A2 => mx_mixer_inst_r375_n122, B => 
                           mx_mixer_inst_r375_n130, C => 
                           mx_mixer_inst_r375_n131, Z => 
                           mx_mixer_inst_r375_n129);
   mx_mixer_inst_r375_U77 : NAN2D1 port map( A1 => mx_mixer_inst_r375_n51, A2 
                           => mx_mixer_inst_r375_n129, Z => 
                           mx_mixer_inst_r375_n127);
   mx_mixer_inst_r375_U76 : NAN2D1 port map( A1 => mx_mixer_inst_r375_n52, A2 
                           => mx_mixer_inst_r375_n129, Z => 
                           mx_mixer_inst_r375_n128);
   mx_mixer_inst_r375_U75 : OAI211D1 port map( A1 => mx_mixer_inst_r375_n121, 
                           A2 => mx_mixer_inst_r375_n119, B => 
                           mx_mixer_inst_r375_n127, C => 
                           mx_mixer_inst_r375_n128, Z => mx_mixer_inst_r375_n13
                           );
   mx_mixer_inst_r375_U74 : NAN2D1 port map( A1 => mixer_in(0), A2 => 
                           mx_mixer_inst_r375_n117, Z => mx_mixer_inst_r375_n48
                           );
   mx_mixer_inst_r375_U73 : EXNOR2D1 port map( A1 => mx_mixer_inst_r375_n117, 
                           A2 => mixer_in(0), Z => mx_mixer_inst_r375_n49);
   mx_mixer_inst_r375_U72 : EXNOR3D1 port map( A1 => mx_mixer_inst_r375_n2, A2 
                           => mixer_in(11), A3 => mixer_in(10), Z => 
                           mx_mixer_inst_N44);
   mx_mixer_inst_r375_U71 : INVD1 port map( A => mixer_in(8), Z => 
                           mx_mixer_inst_r375_n115);
   mx_mixer_inst_r375_U70 : INVD1 port map( A => mixer_in(9), Z => 
                           mx_mixer_inst_r375_n114);
   mx_mixer_inst_r375_U69 : INVD1 port map( A => mixer_in(7), Z => 
                           mx_mixer_inst_r375_n116);
   mx_mixer_inst_r375_U68 : INVD1 port map( A => mixer_in(11), Z => 
                           mx_mixer_inst_r375_n113);
   mx_mixer_inst_r375_U67 : INVD1 port map( A => mixer_in(5), Z => 
                           mx_mixer_inst_r375_n118);
   mx_mixer_inst_r375_U66 : INVD1 port map( A => mixer_in(4), Z => 
                           mx_mixer_inst_r375_n120);
   mx_mixer_inst_r375_U65 : INVD1 port map( A => mixer_in(3), Z => 
                           mx_mixer_inst_r375_n123);
   mx_mixer_inst_r375_U64 : INVD1 port map( A => mixer_in(6), Z => 
                           mx_mixer_inst_r375_n117);
   mx_mixer_inst_r375_U63 : INVD1 port map( A => mixer_in(0), Z => 
                           mx_mixer_inst_r375_n126);
   mx_mixer_inst_r375_U62 : INVD1 port map( A => mixer_in(1), Z => 
                           mx_mixer_inst_r375_n125);
   mx_mixer_inst_r375_U61 : INVD1 port map( A => mixer_in(2), Z => 
                           mx_mixer_inst_r375_n124);
   mx_mixer_inst_r375_U60 : INVD1 port map( A => mx_mixer_inst_r375_n53, Z => 
                           mx_mixer_inst_r375_n122);
   mx_mixer_inst_r375_U59 : INVD1 port map( A => mx_mixer_inst_r375_n51, Z => 
                           mx_mixer_inst_r375_n119);
   mx_mixer_inst_r375_U58 : INVD1 port map( A => mx_mixer_inst_r375_n52, Z => 
                           mx_mixer_inst_r375_n121);
   mx_mixer_inst_r375_U37 : ADHALFDL port map( A => mixer_in(3), B => 
                           mixer_in(4), CO => mx_mixer_inst_r375_n52, S => 
                           mx_mixer_inst_r375_n53);
   mx_mixer_inst_r375_U36 : ADFULD1 port map( A => mixer_in(1), B => 
                           mixer_in(5), CI => mixer_in(4), CO => 
                           mx_mixer_inst_r375_n50, S => mx_mixer_inst_r375_n51)
                           ;
   mx_mixer_inst_r375_U33 : ADFULD1 port map( A => mixer_in(2), B => 
                           mixer_in(5), CI => mx_mixer_inst_r375_n49, CO => 
                           mx_mixer_inst_r375_n46, S => mx_mixer_inst_r375_n47)
                           ;
   mx_mixer_inst_r375_U32 : ADFULD1 port map( A => mixer_in(7), B => 
                           mx_mixer_inst_r375_n125, CI => mixer_in(3), CO => 
                           mx_mixer_inst_r375_n44, S => mx_mixer_inst_r375_n45)
                           ;
   mx_mixer_inst_r375_U31 : ADFULD1 port map( A => mx_mixer_inst_r375_n48, B =>
                           mixer_in(6), CI => mx_mixer_inst_r375_n45, CO => 
                           mx_mixer_inst_r375_n42, S => mx_mixer_inst_r375_n43)
                           ;
   mx_mixer_inst_r375_U30 : ADFULD1 port map( A => mixer_in(8), B => 
                           mx_mixer_inst_r375_n124, CI => mixer_in(4), CO => 
                           mx_mixer_inst_r375_n40, S => mx_mixer_inst_r375_n41)
                           ;
   mx_mixer_inst_r375_U29 : ADFULD1 port map( A => mx_mixer_inst_r375_n44, B =>
                           mixer_in(7), CI => mx_mixer_inst_r375_n41, CO => 
                           mx_mixer_inst_r375_n38, S => mx_mixer_inst_r375_n39)
                           ;
   mx_mixer_inst_r375_U28 : ADFULD1 port map( A => mixer_in(9), B => 
                           mx_mixer_inst_r375_n123, CI => mixer_in(5), CO => 
                           mx_mixer_inst_r375_n36, S => mx_mixer_inst_r375_n37)
                           ;
   mx_mixer_inst_r375_U27 : ADFULD1 port map( A => mx_mixer_inst_r375_n40, B =>
                           mixer_in(8), CI => mx_mixer_inst_r375_n37, CO => 
                           mx_mixer_inst_r375_n34, S => mx_mixer_inst_r375_n35)
                           ;
   mx_mixer_inst_r375_U26 : ADFULD1 port map( A => mixer_in(10), B => 
                           mx_mixer_inst_r375_n120, CI => mixer_in(6), CO => 
                           mx_mixer_inst_r375_n32, S => mx_mixer_inst_r375_n33)
                           ;
   mx_mixer_inst_r375_U25 : ADFULD1 port map( A => mx_mixer_inst_r375_n36, B =>
                           mixer_in(9), CI => mx_mixer_inst_r375_n33, CO => 
                           mx_mixer_inst_r375_n30, S => mx_mixer_inst_r375_n31)
                           ;
   mx_mixer_inst_r375_U24 : ADFULD1 port map( A => mx_mixer_inst_r375_n118, B 
                           => mixer_in(11), CI => mixer_in(10), CO => 
                           mx_mixer_inst_r375_n28, S => mx_mixer_inst_r375_n29)
                           ;
   mx_mixer_inst_r375_U23 : ADFULD1 port map( A => mx_mixer_inst_r375_n32, B =>
                           mixer_in(7), CI => mx_mixer_inst_r375_n29, CO => 
                           mx_mixer_inst_r375_n26, S => mx_mixer_inst_r375_n27)
                           ;
   mx_mixer_inst_r375_U22 : ADFULD1 port map( A => mixer_in(8), B => 
                           mx_mixer_inst_r375_n117, CI => 
                           mx_mixer_inst_r375_n28, CO => mx_mixer_inst_r375_n24
                           , S => mx_mixer_inst_r375_n25);
   mx_mixer_inst_r375_U21 : ADFULD1 port map( A => mx_mixer_inst_r375_n113, B 
                           => mixer_in(7), CI => mixer_in(9), CO => 
                           mx_mixer_inst_r375_n22, S => mx_mixer_inst_r375_n23)
                           ;
   mx_mixer_inst_r375_U20 : ADFULD1 port map( A => mx_mixer_inst_r375_n116, B 
                           => mixer_in(8), CI => mixer_in(10), CO => 
                           mx_mixer_inst_r375_n20, S => mx_mixer_inst_r375_n21)
                           ;
   mx_mixer_inst_r375_U19 : ADFULD1 port map( A => mx_mixer_inst_r375_n115, B 
                           => mx_mixer_inst_r375_n113, CI => 
                           mx_mixer_inst_r375_n114, CO => 
                           mx_mixer_inst_r375_n18, S => mx_mixer_inst_r375_n19)
                           ;
   mx_mixer_inst_r375_U13 : ADFULD1 port map( A => mx_mixer_inst_r375_n47, B =>
                           mx_mixer_inst_r375_n50, CI => mx_mixer_inst_r375_n13
                           , CO => mx_mixer_inst_r375_n12, S => 
                           mx_mixer_inst_N33);
   mx_mixer_inst_r375_U12 : ADFULD1 port map( A => mx_mixer_inst_r375_n43, B =>
                           mx_mixer_inst_r375_n46, CI => mx_mixer_inst_r375_n12
                           , CO => mx_mixer_inst_r375_n11, S => 
                           mx_mixer_inst_N34);
   mx_mixer_inst_r375_U11 : ADFULD1 port map( A => mx_mixer_inst_r375_n39, B =>
                           mx_mixer_inst_r375_n42, CI => mx_mixer_inst_r375_n11
                           , CO => mx_mixer_inst_r375_n10, S => 
                           mx_mixer_inst_N35);
   mx_mixer_inst_r375_U10 : ADFULD1 port map( A => mx_mixer_inst_r375_n35, B =>
                           mx_mixer_inst_r375_n38, CI => mx_mixer_inst_r375_n10
                           , CO => mx_mixer_inst_r375_n9, S => 
                           mx_mixer_inst_N36);
   mx_mixer_inst_r375_U9 : ADFULD1 port map( A => mx_mixer_inst_r375_n31, B => 
                           mx_mixer_inst_r375_n34, CI => mx_mixer_inst_r375_n9,
                           CO => mx_mixer_inst_r375_n8, S => mx_mixer_inst_N37)
                           ;
   mx_mixer_inst_r375_U8 : ADFULD1 port map( A => mx_mixer_inst_r375_n27, B => 
                           mx_mixer_inst_r375_n30, CI => mx_mixer_inst_r375_n8,
                           CO => mx_mixer_inst_r375_n7, S => mx_mixer_inst_N38)
                           ;
   mx_mixer_inst_r375_U7 : ADFULD1 port map( A => mx_mixer_inst_r375_n26, B => 
                           mx_mixer_inst_r375_n25, CI => mx_mixer_inst_r375_n7,
                           CO => mx_mixer_inst_r375_n6, S => mx_mixer_inst_N39)
                           ;
   mx_mixer_inst_r375_U6 : ADFULD1 port map( A => mx_mixer_inst_r375_n24, B => 
                           mx_mixer_inst_r375_n23, CI => mx_mixer_inst_r375_n6,
                           CO => mx_mixer_inst_r375_n5, S => mx_mixer_inst_N40)
                           ;
   mx_mixer_inst_r375_U5 : ADFULD1 port map( A => mx_mixer_inst_r375_n21, B => 
                           mx_mixer_inst_r375_n22, CI => mx_mixer_inst_r375_n5,
                           CO => mx_mixer_inst_r375_n4, S => mx_mixer_inst_N41)
                           ;
   mx_mixer_inst_r375_U4 : ADFULD1 port map( A => mx_mixer_inst_r375_n19, B => 
                           mx_mixer_inst_r375_n20, CI => mx_mixer_inst_r375_n4,
                           CO => mx_mixer_inst_r375_n3, S => mx_mixer_inst_N42)
                           ;
   mx_mixer_inst_r375_U3 : ADFULD1 port map( A => mx_mixer_inst_r375_n18, B => 
                           mixer_in(10), CI => mx_mixer_inst_r375_n3, CO => 
                           mx_mixer_inst_r375_n2, S => mx_mixer_inst_N43);
   mx_mixer_inst_r376_U50 : AOI22D1 port map( A1 => mx_mixer_inst_r376_n52, A2 
                           => mixer_in(0), B1 => mx_mixer_inst_r376_n47, B2 => 
                           mx_mixer_inst_r376_n52, Z => mx_mixer_inst_r376_n104
                           );
   mx_mixer_inst_r376_U49 : OAI21M20D1 port map( A1 => mixer_in(0), A2 => 
                           mx_mixer_inst_r376_n47, B => mx_mixer_inst_r376_n104
                           , Z => mx_mixer_inst_r376_n103);
   mx_mixer_inst_r376_U48 : NAN2D1 port map( A1 => mx_mixer_inst_r376_n50, A2 
                           => mx_mixer_inst_r376_n103, Z => 
                           mx_mixer_inst_r376_n101);
   mx_mixer_inst_r376_U47 : NAN2D1 port map( A1 => mx_mixer_inst_r376_n51, A2 
                           => mx_mixer_inst_r376_n103, Z => 
                           mx_mixer_inst_r376_n102);
   mx_mixer_inst_r376_U46 : OAI211D1 port map( A1 => mx_mixer_inst_r376_n97, A2
                           => mx_mixer_inst_r376_n96, B => 
                           mx_mixer_inst_r376_n101, C => 
                           mx_mixer_inst_r376_n102, Z => 
                           mx_mixer_inst_r376_n100);
   mx_mixer_inst_r376_U45 : NAN2D1 port map( A1 => mx_mixer_inst_r376_n46, A2 
                           => mx_mixer_inst_r376_n100, Z => 
                           mx_mixer_inst_r376_n98);
   mx_mixer_inst_r376_U44 : NAN2D1 port map( A1 => mx_mixer_inst_r376_n49, A2 
                           => mx_mixer_inst_r376_n100, Z => 
                           mx_mixer_inst_r376_n99);
   mx_mixer_inst_r376_U43 : OAI211D1 port map( A1 => mx_mixer_inst_r376_n95, A2
                           => mx_mixer_inst_r376_n94, B => 
                           mx_mixer_inst_r376_n98, C => mx_mixer_inst_r376_n99,
                           Z => mx_mixer_inst_r376_n11);
   mx_mixer_inst_r376_U42 : INVD1 port map( A => mx_mixer_inst_r376_n46, Z => 
                           mx_mixer_inst_r376_n94);
   mx_mixer_inst_r376_U41 : INVD1 port map( A => mx_mixer_inst_r376_n49, Z => 
                           mx_mixer_inst_r376_n95);
   mx_mixer_inst_r376_U40 : INVD1 port map( A => mx_mixer_inst_r376_n50, Z => 
                           mx_mixer_inst_r376_n96);
   mx_mixer_inst_r376_U39 : INVD1 port map( A => mx_mixer_inst_r376_n51, Z => 
                           mx_mixer_inst_r376_n97);
   mx_mixer_inst_r376_U34 : ADHALFDL port map( A => mixer_in(1), B => 
                           mixer_in(3), CO => mx_mixer_inst_r376_n51, S => 
                           mx_mixer_inst_r376_n52);
   mx_mixer_inst_r376_U33 : ADFULD1 port map( A => mixer_in(1), B => 
                           mixer_in(4), CI => mixer_in(2), CO => 
                           mx_mixer_inst_r376_n49, S => mx_mixer_inst_r376_n50)
                           ;
   mx_mixer_inst_r376_U32 : ADHALFDL port map( A => mixer_in(0), B => 
                           mixer_in(2), CO => mx_mixer_inst_r376_n47, S => 
                           mx_mixer_inst_r376_n48);
   mx_mixer_inst_r376_U31 : ADFULD1 port map( A => mixer_in(3), B => 
                           mixer_in(5), CI => mx_mixer_inst_r376_n48, CO => 
                           mx_mixer_inst_r376_n45, S => mx_mixer_inst_r376_n46)
                           ;
   mx_mixer_inst_r376_U30 : ADFULD1 port map( A => mixer_in(1), B => 
                           mixer_in(3), CI => mixer_in(4), CO => 
                           mx_mixer_inst_r376_n43, S => mx_mixer_inst_r376_n44)
                           ;
   mx_mixer_inst_r376_U29 : ADFULD1 port map( A => mx_mixer_inst_r376_n47, B =>
                           mixer_in(6), CI => mx_mixer_inst_r376_n44, CO => 
                           mx_mixer_inst_r376_n41, S => mx_mixer_inst_r376_n42)
                           ;
   mx_mixer_inst_r376_U28 : ADFULD1 port map( A => mixer_in(2), B => 
                           mixer_in(4), CI => mixer_in(5), CO => 
                           mx_mixer_inst_r376_n39, S => mx_mixer_inst_r376_n40)
                           ;
   mx_mixer_inst_r376_U27 : ADFULD1 port map( A => mx_mixer_inst_r376_n43, B =>
                           mixer_in(7), CI => mx_mixer_inst_r376_n40, CO => 
                           mx_mixer_inst_r376_n37, S => mx_mixer_inst_r376_n38)
                           ;
   mx_mixer_inst_r376_U26 : ADFULD1 port map( A => mixer_in(3), B => 
                           mixer_in(5), CI => mixer_in(6), CO => 
                           mx_mixer_inst_r376_n35, S => mx_mixer_inst_r376_n36)
                           ;
   mx_mixer_inst_r376_U25 : ADFULD1 port map( A => mx_mixer_inst_r376_n39, B =>
                           mixer_in(8), CI => mx_mixer_inst_r376_n36, CO => 
                           mx_mixer_inst_r376_n33, S => mx_mixer_inst_r376_n34)
                           ;
   mx_mixer_inst_r376_U24 : ADFULD1 port map( A => mixer_in(4), B => 
                           mixer_in(6), CI => mixer_in(7), CO => 
                           mx_mixer_inst_r376_n31, S => mx_mixer_inst_r376_n32)
                           ;
   mx_mixer_inst_r376_U23 : ADFULD1 port map( A => mx_mixer_inst_r376_n35, B =>
                           mixer_in(9), CI => mx_mixer_inst_r376_n32, CO => 
                           mx_mixer_inst_r376_n29, S => mx_mixer_inst_r376_n30)
                           ;
   mx_mixer_inst_r376_U22 : ADFULD1 port map( A => mixer_in(5), B => 
                           mixer_in(7), CI => mixer_in(8), CO => 
                           mx_mixer_inst_r376_n27, S => mx_mixer_inst_r376_n28)
                           ;
   mx_mixer_inst_r376_U21 : ADFULD1 port map( A => mx_mixer_inst_r376_n31, B =>
                           mixer_in(10), CI => mx_mixer_inst_r376_n28, CO => 
                           mx_mixer_inst_r376_n25, S => mx_mixer_inst_r376_n26)
                           ;
   mx_mixer_inst_r376_U20 : ADFULD1 port map( A => mixer_in(9), B => 
                           mixer_in(11), CI => mixer_in(8), CO => 
                           mx_mixer_inst_r376_n23, S => mx_mixer_inst_r376_n24)
                           ;
   mx_mixer_inst_r376_U19 : ADFULD1 port map( A => mx_mixer_inst_r376_n27, B =>
                           mixer_in(6), CI => mx_mixer_inst_r376_n24, CO => 
                           mx_mixer_inst_r376_n21, S => mx_mixer_inst_r376_n22)
                           ;
   mx_mixer_inst_r376_U18 : ADFULD1 port map( A => mixer_in(10), B => 
                           mixer_in(11), CI => mixer_in(9), CO => 
                           mx_mixer_inst_r376_n19, S => mx_mixer_inst_r376_n20)
                           ;
   mx_mixer_inst_r376_U17 : ADFULD1 port map( A => mx_mixer_inst_r376_n23, B =>
                           mixer_in(7), CI => mx_mixer_inst_r376_n20, CO => 
                           mx_mixer_inst_r376_n17, S => mx_mixer_inst_r376_n18)
                           ;
   mx_mixer_inst_r376_U16 : ADFULD1 port map( A => mixer_in(8), B => 
                           mixer_in(10), CI => mx_mixer_inst_r376_n19, CO => 
                           mx_mixer_inst_r376_n15, S => mx_mixer_inst_r376_n16)
                           ;
   mx_mixer_inst_r376_U11 : ADFULD1 port map( A => mx_mixer_inst_r376_n42, B =>
                           mx_mixer_inst_r376_n45, CI => mx_mixer_inst_r376_n11
                           , CO => mx_mixer_inst_r376_n10, S => 
                           mx_mixer_inst_N45);
   mx_mixer_inst_r376_U10 : ADFULD1 port map( A => mx_mixer_inst_r376_n38, B =>
                           mx_mixer_inst_r376_n41, CI => mx_mixer_inst_r376_n10
                           , CO => mx_mixer_inst_r376_n9, S => 
                           mx_mixer_inst_N46);
   mx_mixer_inst_r376_U9 : ADFULD1 port map( A => mx_mixer_inst_r376_n34, B => 
                           mx_mixer_inst_r376_n37, CI => mx_mixer_inst_r376_n9,
                           CO => mx_mixer_inst_r376_n8, S => mx_mixer_inst_N47)
                           ;
   mx_mixer_inst_r376_U8 : ADFULD1 port map( A => mx_mixer_inst_r376_n30, B => 
                           mx_mixer_inst_r376_n33, CI => mx_mixer_inst_r376_n8,
                           CO => mx_mixer_inst_r376_n7, S => mx_mixer_inst_N48)
                           ;
   mx_mixer_inst_r376_U7 : ADFULD1 port map( A => mx_mixer_inst_r376_n26, B => 
                           mx_mixer_inst_r376_n29, CI => mx_mixer_inst_r376_n7,
                           CO => mx_mixer_inst_r376_n6, S => mx_mixer_inst_N49)
                           ;
   mx_mixer_inst_r376_U6 : ADFULD1 port map( A => mx_mixer_inst_r376_n22, B => 
                           mx_mixer_inst_r376_n25, CI => mx_mixer_inst_r376_n6,
                           CO => mx_mixer_inst_r376_n5, S => mx_mixer_inst_N50)
                           ;
   mx_mixer_inst_r376_U5 : ADFULD1 port map( A => mx_mixer_inst_r376_n18, B => 
                           mx_mixer_inst_r376_n21, CI => mx_mixer_inst_r376_n5,
                           CO => mx_mixer_inst_r376_n4, S => mx_mixer_inst_N51)
                           ;
   mx_mixer_inst_r376_U4 : ADFULD1 port map( A => mx_mixer_inst_r376_n17, B => 
                           mx_mixer_inst_r376_n16, CI => mx_mixer_inst_r376_n4,
                           CO => mx_mixer_inst_r376_n3, S => mx_mixer_inst_N52)
                           ;
   mx_mixer_inst_r376_U3 : ADFULD1 port map( A => mx_mixer_inst_r376_n15, B => 
                           mixer_in(9), CI => mx_mixer_inst_r376_n3, CO => 
                           mx_mixer_inst_r376_n2, S => mx_mixer_inst_N53);
   mx_mixer_inst_r376_U2 : ADFULD1 port map( A => mixer_in(10), B => 
                           mixer_in(11), CI => mx_mixer_inst_r376_n2, CO => 
                           mx_mixer_inst_N55, S => mx_mixer_inst_N54);
   lpf_filter_inst_lpf_i_U94 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair13_15_2_port, A2 => 
                           lpf_filter_inst_lpf_i_p206_1_3, Z => 
                           lpf_filter_inst_lpf_i_p206_1_5);
   lpf_filter_inst_lpf_i_U93 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair13_15_2_port, A2 => 
                           lpf_filter_inst_lpf_i_p206_1_3, Z => 
                           lpf_filter_inst_lpf_i_add_284_carry_3);
   lpf_filter_inst_lpf_i_U92 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_n37, A2 => 
                           lpf_filter_inst_lpf_i_n36, Z => 
                           lpf_filter_inst_lpf_i_t12_13_2);
   lpf_filter_inst_lpf_i_U91 : AND2D1 port map( A1 => lpf_filter_inst_lpf_i_n36
                           , A2 => lpf_filter_inst_lpf_i_n37, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_2_port);
   lpf_filter_inst_lpf_i_U90 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_n38, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_2_port, Z 
                           => lpf_filter_inst_lpf_i_t12_13_3);
   lpf_filter_inst_lpf_i_U89 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_2_port, 
                           A2 => lpf_filter_inst_lpf_i_n38, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_3_port);
   lpf_filter_inst_lpf_i_U88 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t11_14_0_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_168_port, Z => 
                           lpf_filter_inst_lpf_i_p232_2_1);
   lpf_filter_inst_lpf_i_U87 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t11_14_0_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_168_port, Z => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_2);
   lpf_filter_inst_lpf_i_U86 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_n50, A2 => 
                           lpf_filter_inst_lpf_i_n49, Z => 
                           lpf_filter_inst_lpf_i_n157);
   lpf_filter_inst_lpf_i_U85 : AND2D1 port map( A1 => lpf_filter_inst_lpf_i_n49
                           , A2 => lpf_filter_inst_lpf_i_n50, Z => 
                           lpf_filter_inst_lpf_i_sub_280_carry_2_port);
   lpf_filter_inst_lpf_i_U84 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_n51, A2 => 
                           lpf_filter_inst_lpf_i_sub_280_carry_2_port, Z => 
                           lpf_filter_inst_lpf_i_p141_1_2_port);
   lpf_filter_inst_lpf_i_U83 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_280_carry_2_port, A2 => 
                           lpf_filter_inst_lpf_i_n51, Z => 
                           lpf_filter_inst_lpf_i_sub_280_carry_3_port);
   lpf_filter_inst_lpf_i_U82 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_n52, A2 => 
                           lpf_filter_inst_lpf_i_sub_280_carry_3_port, Z => 
                           lpf_filter_inst_lpf_i_p141_1_3_port);
   lpf_filter_inst_lpf_i_U81 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_280_carry_3_port, A2 => 
                           lpf_filter_inst_lpf_i_n52, Z => 
                           lpf_filter_inst_lpf_i_sub_280_carry_4_port);
   lpf_filter_inst_lpf_i_U80 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_n53, A2 => 
                           lpf_filter_inst_lpf_i_sub_280_carry_4_port, Z => 
                           lpf_filter_inst_lpf_i_p141_1_4_port);
   lpf_filter_inst_lpf_i_U79 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_280_carry_4_port, A2 => 
                           lpf_filter_inst_lpf_i_n53, Z => 
                           lpf_filter_inst_lpf_i_sub_280_carry_5_port);
   lpf_filter_inst_lpf_i_U78 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_n54, A2 => 
                           lpf_filter_inst_lpf_i_sub_280_carry_5_port, Z => 
                           lpf_filter_inst_lpf_i_p141_1_5_port);
   lpf_filter_inst_lpf_i_U77 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_280_carry_5_port, A2 => 
                           lpf_filter_inst_lpf_i_n54, Z => 
                           lpf_filter_inst_lpf_i_sub_280_carry_6_port);
   lpf_filter_inst_lpf_i_U76 : TIELO port map( Z => 
                           lpf_filter_inst_lpf_i_net5306);
   lpf_filter_inst_lpf_i_U75 : INVD1 port map( A => rstn, Z => 
                           lpf_filter_inst_lpf_i_n3);
   lpf_filter_inst_lpf_i_U74 : BUFD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_12_port, Z => 
                           lpf_filter_inst_lpf_i_n1);
   lpf_filter_inst_lpf_i_U73 : BUFD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_178_port, Z => 
                           lpf_filter_inst_lpf_i_p232_2_17);
   lpf_filter_inst_lpf_i_U72 : INVD1 port map( A => lpf_filter_inst_lpf_i_n3, Z
                           => lpf_filter_inst_lpf_i_n2);
   lpf_filter_inst_lpf_i_U71 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_2_port, Z => 
                           lpf_filter_inst_lpf_i_n38);
   lpf_filter_inst_lpf_i_U70 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_3, Z => 
                           lpf_filter_inst_lpf_i_n36);
   lpf_filter_inst_lpf_i_U69 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_5_port, Z => 
                           lpf_filter_inst_lpf_i_n54);
   lpf_filter_inst_lpf_i_U68 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_4_port, Z => 
                           lpf_filter_inst_lpf_i_n53);
   lpf_filter_inst_lpf_i_U67 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_3_port, Z => 
                           lpf_filter_inst_lpf_i_n52);
   lpf_filter_inst_lpf_i_U66 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_2_port, Z => 
                           lpf_filter_inst_lpf_i_n51);
   lpf_filter_inst_lpf_i_U65 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_4, Z => 
                           lpf_filter_inst_lpf_i_n37);
   lpf_filter_inst_lpf_i_U64 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_1_port, Z => 
                           lpf_filter_inst_lpf_i_n50);
   lpf_filter_inst_lpf_i_U63 : INVD1 port map( A => lpf_filter_inst_lpf_i_n117,
                           Z => lpf_filter_inst_lpf_i_n49);
   lpf_filter_inst_lpf_i_U62 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_11_port, Z => 
                           lpf_filter_inst_lpf_i_n47);
   lpf_filter_inst_lpf_i_U61 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_10_port, Z => 
                           lpf_filter_inst_lpf_i_n46);
   lpf_filter_inst_lpf_i_U60 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_9_port, Z => 
                           lpf_filter_inst_lpf_i_n45);
   lpf_filter_inst_lpf_i_U59 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_8_port, Z => 
                           lpf_filter_inst_lpf_i_n44);
   lpf_filter_inst_lpf_i_U58 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_7_port, Z => 
                           lpf_filter_inst_lpf_i_n43);
   lpf_filter_inst_lpf_i_U57 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_6_port, Z => 
                           lpf_filter_inst_lpf_i_n42);
   lpf_filter_inst_lpf_i_U56 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_5_port, Z => 
                           lpf_filter_inst_lpf_i_n41);
   lpf_filter_inst_lpf_i_U55 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_11_port, Z => 
                           lpf_filter_inst_lpf_i_n60);
   lpf_filter_inst_lpf_i_U54 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_10_port, Z => 
                           lpf_filter_inst_lpf_i_n59);
   lpf_filter_inst_lpf_i_U53 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_9_port, Z => 
                           lpf_filter_inst_lpf_i_n58);
   lpf_filter_inst_lpf_i_U52 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_8_port, Z => 
                           lpf_filter_inst_lpf_i_n57);
   lpf_filter_inst_lpf_i_U51 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_4_port, Z => 
                           lpf_filter_inst_lpf_i_n40);
   lpf_filter_inst_lpf_i_U50 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_7_port, Z => 
                           lpf_filter_inst_lpf_i_n56);
   lpf_filter_inst_lpf_i_U49 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_3_port, Z => 
                           lpf_filter_inst_lpf_i_n39);
   lpf_filter_inst_lpf_i_U48 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_6_port, Z => 
                           lpf_filter_inst_lpf_i_n55);
   lpf_filter_inst_lpf_i_U47 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_2_15_port, Z => 
                           lpf_filter_inst_lpf_i_n48);
   lpf_filter_inst_lpf_i_U46 : INVD1 port map( A => lpf_filter_inst_lpf_i_n1, Z
                           => lpf_filter_inst_lpf_i_n61);
   lpf_filter_inst_lpf_i_U45 : INVD1 port map( A => lpf_filter_inst_lpf_i_n2, Z
                           => lpf_filter_inst_lpf_i_n35);
   lpf_filter_inst_lpf_i_U44 : INVD1 port map( A => lpf_filter_inst_lpf_i_n2, Z
                           => lpf_filter_inst_lpf_i_n34);
   lpf_filter_inst_lpf_i_U43 : INVD1 port map( A => lpf_filter_inst_lpf_i_n2, Z
                           => lpf_filter_inst_lpf_i_n33);
   lpf_filter_inst_lpf_i_U42 : INVD1 port map( A => lpf_filter_inst_lpf_i_n2, Z
                           => lpf_filter_inst_lpf_i_n32);
   lpf_filter_inst_lpf_i_U41 : INVD1 port map( A => lpf_filter_inst_lpf_i_n2, Z
                           => lpf_filter_inst_lpf_i_n31);
   lpf_filter_inst_lpf_i_U40 : INVD1 port map( A => lpf_filter_inst_lpf_i_n2, Z
                           => lpf_filter_inst_lpf_i_n30);
   lpf_filter_inst_lpf_i_U39 : OAI21M20D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_12_port, 
                           A2 => lpf_filter_inst_lpf_i_n68, B => 
                           lpf_filter_inst_lpf_i_n69, Z => filter_out_i_0_port)
                           ;
   lpf_filter_inst_lpf_i_U38 : OAI21M20D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_13_port, 
                           A2 => lpf_filter_inst_lpf_i_n68, B => 
                           lpf_filter_inst_lpf_i_n69, Z => filter_out_i_1_port)
                           ;
   lpf_filter_inst_lpf_i_U37 : NAN4D1 port map( A1 => filter_out_i_4_port, A2 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_22_port, 
                           A3 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_21_port, 
                           A4 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_20_port, Z 
                           => lpf_filter_inst_lpf_i_n71);
   lpf_filter_inst_lpf_i_U36 : OAI21M20D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_15_port, 
                           A2 => lpf_filter_inst_lpf_i_n68, B => 
                           lpf_filter_inst_lpf_i_n69, Z => filter_out_i_3_port)
                           ;
   lpf_filter_inst_lpf_i_U35 : OAI21M20D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_14_port, 
                           A2 => lpf_filter_inst_lpf_i_n68, B => 
                           lpf_filter_inst_lpf_i_n69, Z => filter_out_i_2_port)
                           ;
   lpf_filter_inst_lpf_i_U34 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_sub_280_carry_18_port, Z => 
                           lpf_filter_inst_lpf_i_p141_1_19_port);
   lpf_filter_inst_lpf_i_U33 : NAN4D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_19_port, 
                           A2 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_18_port, 
                           A3 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_17_port, 
                           A4 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_16_port, Z 
                           => lpf_filter_inst_lpf_i_n70);
   lpf_filter_inst_lpf_i_U32 : INVD1 port map( A => lpf_filter_inst_lpf_i_n30, 
                           Z => lpf_filter_inst_lpf_i_n29);
   lpf_filter_inst_lpf_i_U31 : INVD1 port map( A => lpf_filter_inst_lpf_i_n30, 
                           Z => lpf_filter_inst_lpf_i_n4);
   lpf_filter_inst_lpf_i_U30 : INVD1 port map( A => lpf_filter_inst_lpf_i_n3, Z
                           => lpf_filter_inst_lpf_i_n5);
   lpf_filter_inst_lpf_i_U29 : INVD1 port map( A => lpf_filter_inst_lpf_i_n31, 
                           Z => lpf_filter_inst_lpf_i_n6);
   lpf_filter_inst_lpf_i_U28 : INVD1 port map( A => lpf_filter_inst_lpf_i_n35, 
                           Z => lpf_filter_inst_lpf_i_n7);
   lpf_filter_inst_lpf_i_U27 : INVD1 port map( A => lpf_filter_inst_lpf_i_n3, Z
                           => lpf_filter_inst_lpf_i_n8);
   lpf_filter_inst_lpf_i_U26 : INVD1 port map( A => lpf_filter_inst_lpf_i_n35, 
                           Z => lpf_filter_inst_lpf_i_n9);
   lpf_filter_inst_lpf_i_U25 : INVD1 port map( A => lpf_filter_inst_lpf_i_n35, 
                           Z => lpf_filter_inst_lpf_i_n10);
   lpf_filter_inst_lpf_i_U24 : INVD1 port map( A => lpf_filter_inst_lpf_i_n35, 
                           Z => lpf_filter_inst_lpf_i_n11);
   lpf_filter_inst_lpf_i_U23 : INVD1 port map( A => lpf_filter_inst_lpf_i_n34, 
                           Z => lpf_filter_inst_lpf_i_n12);
   lpf_filter_inst_lpf_i_U22 : INVD1 port map( A => lpf_filter_inst_lpf_i_n33, 
                           Z => lpf_filter_inst_lpf_i_n13);
   lpf_filter_inst_lpf_i_U21 : INVD1 port map( A => lpf_filter_inst_lpf_i_n32, 
                           Z => lpf_filter_inst_lpf_i_n14);
   lpf_filter_inst_lpf_i_U20 : INVD1 port map( A => lpf_filter_inst_lpf_i_n34, 
                           Z => lpf_filter_inst_lpf_i_n15);
   lpf_filter_inst_lpf_i_U15 : INVD1 port map( A => lpf_filter_inst_lpf_i_n34, 
                           Z => lpf_filter_inst_lpf_i_n16);
   lpf_filter_inst_lpf_i_U14 : INVD1 port map( A => lpf_filter_inst_lpf_i_n34, 
                           Z => lpf_filter_inst_lpf_i_n17);
   lpf_filter_inst_lpf_i_U13 : INVD1 port map( A => lpf_filter_inst_lpf_i_n33, 
                           Z => lpf_filter_inst_lpf_i_n18);
   lpf_filter_inst_lpf_i_U12 : INVD1 port map( A => lpf_filter_inst_lpf_i_n33, 
                           Z => lpf_filter_inst_lpf_i_n19);
   lpf_filter_inst_lpf_i_U11 : INVD1 port map( A => lpf_filter_inst_lpf_i_n33, 
                           Z => lpf_filter_inst_lpf_i_n20);
   lpf_filter_inst_lpf_i_U10 : INVD1 port map( A => lpf_filter_inst_lpf_i_n32, 
                           Z => lpf_filter_inst_lpf_i_n21);
   lpf_filter_inst_lpf_i_U9 : INVD1 port map( A => lpf_filter_inst_lpf_i_n32, Z
                           => lpf_filter_inst_lpf_i_n22);
   lpf_filter_inst_lpf_i_U8 : INVD1 port map( A => lpf_filter_inst_lpf_i_n32, Z
                           => lpf_filter_inst_lpf_i_n23);
   lpf_filter_inst_lpf_i_U7 : INVD1 port map( A => lpf_filter_inst_lpf_i_n31, Z
                           => lpf_filter_inst_lpf_i_n24);
   lpf_filter_inst_lpf_i_U6 : INVD1 port map( A => lpf_filter_inst_lpf_i_n31, Z
                           => lpf_filter_inst_lpf_i_n25);
   lpf_filter_inst_lpf_i_U5 : INVD1 port map( A => lpf_filter_inst_lpf_i_n31, Z
                           => lpf_filter_inst_lpf_i_n26);
   lpf_filter_inst_lpf_i_U4 : INVD1 port map( A => lpf_filter_inst_lpf_i_n30, Z
                           => lpf_filter_inst_lpf_i_n27);
   lpf_filter_inst_lpf_i_U3 : INVD1 port map( A => lpf_filter_inst_lpf_i_n30, Z
                           => lpf_filter_inst_lpf_i_n28);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_36_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_24_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_37_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_25_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_38_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_26_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_39_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_27_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_40_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_28_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_41_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_29_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_42_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_30_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_43_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_31_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_44_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_32_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_45_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_33_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_46_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_34_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_25_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_47_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_35_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_84_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_72_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_85_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_73_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_86_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_74_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_87_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_75_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_88_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_76_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_89_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_77_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_90_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_78_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_91_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_79_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_92_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_80_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_93_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_81_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_94_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_82_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_21_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_95_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_83_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_132_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_120_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_133_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_121_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_134_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_122_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_135_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_123_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_136_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_124_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_137_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_125_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_138_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_126_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_139_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_127_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_140_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_128_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_141_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_129_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_142_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_130_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_17_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_143_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_131_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_227_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_215_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_228_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_216_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_229_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_217_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_230_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_218_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_231_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_219_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_232_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_220_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_233_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_221_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_234_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_222_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_235_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_223_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_236_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_224_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_237_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_225_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_9_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_238_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_226_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_275_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_263_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_276_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_264_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_277_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_265_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_278_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_266_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_279_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_267_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_280_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_268_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_281_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_269_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_282_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_270_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_283_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_271_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_284_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_272_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_285_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_273_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_5_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_286_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_274_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_323_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_311_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_324_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_312_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_325_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_313_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_326_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_314_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_327_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_315_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_328_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_316_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_329_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_317_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_330_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_318_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_331_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_319_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_332_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_320_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_333_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_321_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_1_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_334_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_322_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_190_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_178_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_179_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_t11_14_0_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_181_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_169_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_182_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_170_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_183_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_171_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_184_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_172_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_185_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_173_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_186_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_174_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_187_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_175_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_188_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_176_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_189_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_177_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_13_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_180_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_168_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_202_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_190_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_214_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_202_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_226_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_214_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_250_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_238_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_262_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_250_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_274_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_262_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_298_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_286_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_310_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_298_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_322_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_310_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_11 : DFFRPQ1 port map( D => 
                           mixer_out_i_11_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_334_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_35_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_23_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_59_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_47_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_71_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_59_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_83_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_71_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_107_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_95_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_119_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_107_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_131_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_119_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_155_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_143_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_167_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_155_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_p232_2_17, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n16, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_167_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_24_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_12_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_48_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n27, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_36_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_60_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_48_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_72_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_60_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_96_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_84_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_108_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_96_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_120_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_108_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_144_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_132_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_156_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_144_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_t11_14_0_port, CK => clk, RB 
                           => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_156_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_192_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_180_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_193_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_181_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_194_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_182_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_195_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_183_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_196_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_184_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_197_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_185_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_198_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_186_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_199_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_187_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_200_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_188_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_201_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_189_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_204_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_192_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_205_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_193_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_206_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_194_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_207_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_195_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_208_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_196_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_209_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_197_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_210_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_198_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_211_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_199_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_212_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_200_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_213_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_201_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_216_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_204_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_217_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_205_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_218_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_206_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_219_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_207_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_220_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_208_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_221_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_209_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_222_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_210_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_223_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_211_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_224_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_212_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_225_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n13, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_213_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_240_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_228_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_241_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_229_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_242_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_230_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_243_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_231_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_244_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_232_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_245_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_233_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_246_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_234_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_247_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_235_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_248_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_236_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_249_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_237_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_252_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_240_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_253_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_241_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_254_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_242_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_255_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_243_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_256_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_244_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_257_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_245_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_258_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_246_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_259_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_247_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_260_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_248_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_261_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_249_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_264_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_252_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_265_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_253_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_266_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_254_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_267_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_255_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_268_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_256_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_269_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_257_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_270_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_258_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_271_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_259_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_272_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_260_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_273_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n9, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_261_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_288_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_276_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_289_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_277_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_290_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_278_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_291_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_279_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_292_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_280_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_293_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_281_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_294_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_282_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_295_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_283_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_296_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_284_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_297_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_285_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_300_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_288_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_301_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_289_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_302_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_290_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_303_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_291_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_304_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_292_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_305_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_293_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_306_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_294_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_307_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_295_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_308_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_296_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_309_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_297_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_312_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_300_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_313_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_301_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_314_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_302_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_315_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_303_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_316_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_304_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_317_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_305_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_318_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_306_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_319_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_307_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_320_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_308_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_321_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n5, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_309_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_1 : DFFRPQ1 port map( D => 
                           mixer_out_i_1_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_324_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_2 : DFFRPQ1 port map( D => 
                           mixer_out_i_2_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_325_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_3 : DFFRPQ1 port map( D => 
                           mixer_out_i_3_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_326_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_4 : DFFRPQ1 port map( D => 
                           mixer_out_i_4_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_327_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_5 : DFFRPQ1 port map( D => 
                           mixer_out_i_5_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_328_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_6 : DFFRPQ1 port map( D => 
                           mixer_out_i_6_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_329_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_7 : DFFRPQ1 port map( D => 
                           mixer_out_i_7_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_330_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_8 : DFFRPQ1 port map( D => 
                           mixer_out_i_8_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_331_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_9 : DFFRPQ1 port map( D => 
                           mixer_out_i_9_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_332_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_10 : DFFRPQ1 port map( D => 
                           mixer_out_i_10_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_333_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_25_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_13_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_26_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_14_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_27_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_15_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_28_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_16_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_29_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_17_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_30_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_18_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_31_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_19_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_32_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_20_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_33_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_21_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_26_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_34_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_22_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_49_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_37_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_50_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_38_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_51_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_39_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_52_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_40_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_53_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_41_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_54_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_42_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_55_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_43_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_56_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_44_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_57_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_45_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_24_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_58_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_46_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_61_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n26, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_49_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_62_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_50_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_63_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_51_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_64_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_52_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_65_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_53_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_66_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_54_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_67_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_55_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_68_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_56_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_69_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_57_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_23_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_70_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_58_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_73_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_61_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_74_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n25, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_62_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_75_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_63_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_76_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_64_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_77_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_65_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_78_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_66_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_79_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_67_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_80_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_68_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_81_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_69_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_22_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_82_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n24, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_70_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_97_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_85_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_98_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_86_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_99_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_87_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_100_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n23, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_88_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_101_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_89_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_102_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_90_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_103_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_91_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_104_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_92_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_105_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_93_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_20_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_106_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_94_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_109_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_97_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_110_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_98_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_111_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_99_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_112_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_100_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_113_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n22, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_101_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_114_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_102_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_115_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_103_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_116_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_104_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_117_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_105_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_19_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_118_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_106_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_121_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_109_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_122_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_110_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_123_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_111_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_124_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_112_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_125_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_113_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_126_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n21, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_114_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_127_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_115_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_128_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_116_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_129_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_117_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_18_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_130_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n20, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_118_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_145_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_133_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_146_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_134_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_147_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_135_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_148_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_136_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_149_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_137_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_150_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_138_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_151_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_139_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_152_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n19, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_140_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_153_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_141_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_16_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_154_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_142_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_157_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_145_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_158_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_146_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_159_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_147_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_160_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_148_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_161_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_149_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_162_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_150_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_163_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_151_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_164_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_152_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_165_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n18, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_153_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_15_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_166_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_154_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_168_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_157_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_169_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_158_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_170_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_159_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_171_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_160_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_172_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_161_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_173_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_162_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_174_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_163_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_175_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_164_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_176_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_165_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_14_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_177_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n17, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_166_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_12_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_191_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_179_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_11_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_203_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n15, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_191_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_10_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_215_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n14, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_203_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_8_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_239_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n12, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_227_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_7_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_251_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n11, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_239_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_6_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_263_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n10, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_251_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_4_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_287_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n8, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_275_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_3_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_299_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n7, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_287_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_2_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_311_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n6, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_299_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_0_0 : DFFRPQ1 port map( D => 
                           mixer_out_i_0_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_i_n4, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_323_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_23_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n28, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_11_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_12_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_0_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_13_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_1_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_14_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_2_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_15_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_3_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_16_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_4_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_17_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_5_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_18_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_6_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_19_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_7_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_20_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_8_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_21_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_9_port);
   lpf_filter_inst_lpf_i_arx_input_reg_reg_27_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_i_arx_input_reg_22_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_i_n29, Q => 
                           lpf_filter_inst_lpf_i_arx_input_reg_10_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_20 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_19, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_20_port, 
                           CO => lpf_filter_inst_lpf_i_n_1421, S => 
                           lpf_filter_inst_lpf_i_p206_3_20_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_19, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_20_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_19_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_18, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_19_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_18_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_17, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_17_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_16, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_16_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_15, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_15_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_14, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_14_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_13, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_13_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_12, B => 
                           lpf_filter_inst_lpf_i_n48, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_12_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_11, B => 
                           lpf_filter_inst_lpf_i_n47, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_11_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_10, B => 
                           lpf_filter_inst_lpf_i_n46, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_10_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_9, B => 
                           lpf_filter_inst_lpf_i_n45, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_9_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_8, B => 
                           lpf_filter_inst_lpf_i_n44, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_8_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_7, B => 
                           lpf_filter_inst_lpf_i_n43, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_7_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_6, B => 
                           lpf_filter_inst_lpf_i_n42, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_6_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_5, B => 
                           lpf_filter_inst_lpf_i_n41, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_5_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_4, B => 
                           lpf_filter_inst_lpf_i_n40, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_4_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_285_U2_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_3, B => 
                           lpf_filter_inst_lpf_i_n39, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_285_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_p206_3_3_port);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_17, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_177_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_11, 
                           CO => lpf_filter_inst_lpf_i_p232_2_12, S => 
                           lpf_filter_inst_lpf_i_p232_2_11);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_177_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_176_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_10, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_11, S
                           => lpf_filter_inst_lpf_i_p232_2_10);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_176_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_175_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_9, CO
                           => lpf_filter_inst_lpf_i_add_1_root_add_286_carry_10
                           , S => lpf_filter_inst_lpf_i_p232_2_9);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_175_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_174_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_8, CO
                           => lpf_filter_inst_lpf_i_add_1_root_add_286_carry_9,
                           S => lpf_filter_inst_lpf_i_p232_2_8);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_174_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_173_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_7, CO
                           => lpf_filter_inst_lpf_i_add_1_root_add_286_carry_8,
                           S => lpf_filter_inst_lpf_i_p232_2_7);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_173_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_172_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_6, CO
                           => lpf_filter_inst_lpf_i_add_1_root_add_286_carry_7,
                           S => lpf_filter_inst_lpf_i_p232_2_6);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_172_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_171_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_5, CO
                           => lpf_filter_inst_lpf_i_add_1_root_add_286_carry_6,
                           S => lpf_filter_inst_lpf_i_p232_2_5);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_171_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_170_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_4, CO
                           => lpf_filter_inst_lpf_i_add_1_root_add_286_carry_5,
                           S => lpf_filter_inst_lpf_i_p232_2_4);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_170_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_169_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_3, CO
                           => lpf_filter_inst_lpf_i_add_1_root_add_286_carry_4,
                           S => lpf_filter_inst_lpf_i_p232_2_3);
   lpf_filter_inst_lpf_i_add_1_root_add_286_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_169_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_168_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_286_carry_2, CO
                           => lpf_filter_inst_lpf_i_add_1_root_add_286_carry_3,
                           S => lpf_filter_inst_lpf_i_p232_2_2);
   lpf_filter_inst_lpf_i_sub_280_U2_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_11_port, B => 
                           lpf_filter_inst_lpf_i_n61, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_17_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_18_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_17_port);
   lpf_filter_inst_lpf_i_sub_280_U2_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_10_port, B => 
                           lpf_filter_inst_lpf_i_n61, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_16_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_17_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_16_port);
   lpf_filter_inst_lpf_i_sub_280_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_9_port, B => 
                           lpf_filter_inst_lpf_i_n61, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_15_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_16_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_15_port);
   lpf_filter_inst_lpf_i_sub_280_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_8_port, B => 
                           lpf_filter_inst_lpf_i_n61, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_14_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_15_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_14_port);
   lpf_filter_inst_lpf_i_sub_280_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_7_port, B => 
                           lpf_filter_inst_lpf_i_n61, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_13_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_14_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_13_port);
   lpf_filter_inst_lpf_i_sub_280_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_6_port, B => 
                           lpf_filter_inst_lpf_i_n61, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_12_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_13_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_12_port);
   lpf_filter_inst_lpf_i_sub_280_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_5_port, B => 
                           lpf_filter_inst_lpf_i_n60, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_11_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_12_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_11_port);
   lpf_filter_inst_lpf_i_sub_280_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_4_port, B => 
                           lpf_filter_inst_lpf_i_n59, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_10_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_11_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_10_port);
   lpf_filter_inst_lpf_i_sub_280_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_3_port, B => 
                           lpf_filter_inst_lpf_i_n58, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_9_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_10_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_9_port);
   lpf_filter_inst_lpf_i_sub_280_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_2_port, B => 
                           lpf_filter_inst_lpf_i_n57, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_8_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_9_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_8_port);
   lpf_filter_inst_lpf_i_sub_280_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_1_port, B => 
                           lpf_filter_inst_lpf_i_n56, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_7_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_8_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_7_port);
   lpf_filter_inst_lpf_i_sub_280_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n117, B => 
                           lpf_filter_inst_lpf_i_n55, CI => 
                           lpf_filter_inst_lpf_i_sub_280_carry_6_port, CO => 
                           lpf_filter_inst_lpf_i_sub_280_carry_7_port, S => 
                           lpf_filter_inst_lpf_i_p141_1_6_port);
   lpf_filter_inst_lpf_i_add_284_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_11_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_15_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_13, CO => 
                           lpf_filter_inst_lpf_i_p206_2_14_port, S => 
                           lpf_filter_inst_lpf_i_p206_2_13_port);
   lpf_filter_inst_lpf_i_add_284_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_10_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_15_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_12, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_13, S => 
                           lpf_filter_inst_lpf_i_p206_2_12_port);
   lpf_filter_inst_lpf_i_add_284_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_9_port, B => 
                           lpf_filter_inst_lpf_i_pair13_15_11_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_11, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_12, S => 
                           lpf_filter_inst_lpf_i_p206_2_11_port);
   lpf_filter_inst_lpf_i_add_284_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_8_port, B => 
                           lpf_filter_inst_lpf_i_pair13_15_10_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_10, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_11, S => 
                           lpf_filter_inst_lpf_i_p206_2_10_port);
   lpf_filter_inst_lpf_i_add_284_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_7_port, B => 
                           lpf_filter_inst_lpf_i_pair13_15_9_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_9, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_10, S => 
                           lpf_filter_inst_lpf_i_p206_2_9_port);
   lpf_filter_inst_lpf_i_add_284_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_6_port, B => 
                           lpf_filter_inst_lpf_i_pair13_15_8_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_8, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_9, S => 
                           lpf_filter_inst_lpf_i_p206_2_8_port);
   lpf_filter_inst_lpf_i_add_284_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_5_port, B => 
                           lpf_filter_inst_lpf_i_pair13_15_7_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_7, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_8, S => 
                           lpf_filter_inst_lpf_i_p206_2_7_port);
   lpf_filter_inst_lpf_i_add_284_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_4_port, B => 
                           lpf_filter_inst_lpf_i_pair13_15_6_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_6, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_7, S => 
                           lpf_filter_inst_lpf_i_p206_2_6_port);
   lpf_filter_inst_lpf_i_add_284_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_3_port, B => 
                           lpf_filter_inst_lpf_i_pair13_15_5_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_5, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_6, S => 
                           lpf_filter_inst_lpf_i_p206_2_5_port);
   lpf_filter_inst_lpf_i_add_284_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_2_port, B => 
                           lpf_filter_inst_lpf_i_pair13_15_4_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_4, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_5, S => 
                           lpf_filter_inst_lpf_i_p206_2_4_port);
   lpf_filter_inst_lpf_i_add_284_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_4, B => 
                           lpf_filter_inst_lpf_i_pair13_15_3_port, CI => 
                           lpf_filter_inst_lpf_i_add_284_carry_3, CO => 
                           lpf_filter_inst_lpf_i_add_284_carry_4, S => 
                           lpf_filter_inst_lpf_i_p206_2_3_port);
   lpf_filter_inst_lpf_i_U19 : OR4D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_20_port, 
                           A2 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_21_port, 
                           A3 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_22_port, 
                           A4 => filter_out_i_4_port, Z => 
                           lpf_filter_inst_lpf_i_n72);
   lpf_filter_inst_lpf_i_U18 : OR4D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_16_port, 
                           A2 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_17_port, 
                           A3 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_18_port, 
                           A4 => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_19_port, Z 
                           => lpf_filter_inst_lpf_i_n73);
   lpf_filter_inst_lpf_i_U17 : OAI22D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_n70, A2 => 
                           lpf_filter_inst_lpf_i_n71, B1 => 
                           lpf_filter_inst_lpf_i_n72, B2 => 
                           lpf_filter_inst_lpf_i_n73, Z => 
                           lpf_filter_inst_lpf_i_n68);
   lpf_filter_inst_lpf_i_U16 : OR2D1 port map( A1 => lpf_filter_inst_lpf_i_n68,
                           A2 => filter_out_i_4_port, Z => 
                           lpf_filter_inst_lpf_i_n69);
   lpf_filter_inst_lpf_i_add_273_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_156_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_179_port, Z => 
                           lpf_filter_inst_lpf_i_p206_1_3);
   lpf_filter_inst_lpf_i_add_273_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_156_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_179_port, Z => 
                           lpf_filter_inst_lpf_i_add_273_n1);
   lpf_filter_inst_lpf_i_add_273_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_180_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_157_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_n1, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_2_port, S => 
                           lpf_filter_inst_lpf_i_p206_1_4);
   lpf_filter_inst_lpf_i_add_273_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_181_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_158_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_2_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_3_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_2_port);
   lpf_filter_inst_lpf_i_add_273_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_182_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_159_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_3_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_4_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_3_port);
   lpf_filter_inst_lpf_i_add_273_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_183_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_160_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_4_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_5_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_4_port);
   lpf_filter_inst_lpf_i_add_273_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_184_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_161_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_5_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_6_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_5_port);
   lpf_filter_inst_lpf_i_add_273_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_185_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_162_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_6_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_7_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_6_port);
   lpf_filter_inst_lpf_i_add_273_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_186_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_163_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_7_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_8_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_7_port);
   lpf_filter_inst_lpf_i_add_273_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_187_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_164_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_8_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_9_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_8_port);
   lpf_filter_inst_lpf_i_add_273_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_188_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_165_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_9_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_10_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_9_port);
   lpf_filter_inst_lpf_i_add_273_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_189_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_166_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_10_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_11_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_10_port);
   lpf_filter_inst_lpf_i_add_273_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_190_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_167_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_11_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_carry_12_port, S => 
                           lpf_filter_inst_lpf_i_pair13_15_11_port);
   lpf_filter_inst_lpf_i_add_273_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_190_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_167_port, CI => 
                           lpf_filter_inst_lpf_i_add_273_carry_12_port, CO => 
                           lpf_filter_inst_lpf_i_add_273_n_1308, S => 
                           lpf_filter_inst_lpf_i_p206_2_15_port);
   lpf_filter_inst_lpf_i_add_272_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_144_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_191_port, Z => 
                           lpf_filter_inst_lpf_i_n117);
   lpf_filter_inst_lpf_i_add_272_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_144_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_191_port, Z => 
                           lpf_filter_inst_lpf_i_add_272_n1);
   lpf_filter_inst_lpf_i_add_272_U1_12 : EXOR3D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_202_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_155_port, A3 => 
                           lpf_filter_inst_lpf_i_add_272_carry_12_port, Z => 
                           lpf_filter_inst_lpf_i_pair12_16_12_port);
   lpf_filter_inst_lpf_i_add_272_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_192_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_145_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_n1, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_2_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_1_port);
   lpf_filter_inst_lpf_i_add_272_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_193_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_146_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_2_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_3_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_2_port);
   lpf_filter_inst_lpf_i_add_272_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_194_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_147_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_3_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_4_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_3_port);
   lpf_filter_inst_lpf_i_add_272_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_195_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_148_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_4_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_5_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_4_port);
   lpf_filter_inst_lpf_i_add_272_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_196_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_149_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_5_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_6_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_5_port);
   lpf_filter_inst_lpf_i_add_272_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_197_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_150_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_6_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_7_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_6_port);
   lpf_filter_inst_lpf_i_add_272_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_198_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_151_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_7_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_8_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_7_port);
   lpf_filter_inst_lpf_i_add_272_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_199_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_152_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_8_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_9_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_8_port);
   lpf_filter_inst_lpf_i_add_272_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_200_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_153_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_9_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_10_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_9_port);
   lpf_filter_inst_lpf_i_add_272_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_201_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_154_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_10_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_11_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_10_port);
   lpf_filter_inst_lpf_i_add_272_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_202_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_155_port, CI => 
                           lpf_filter_inst_lpf_i_add_272_carry_11_port, CO => 
                           lpf_filter_inst_lpf_i_add_272_carry_12_port, S => 
                           lpf_filter_inst_lpf_i_pair12_16_11_port);
   lpf_filter_inst_lpf_i_add_271_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_132_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_203_port, Z => 
                           lpf_filter_inst_lpf_i_n74);
   lpf_filter_inst_lpf_i_add_271_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_132_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_203_port, Z => 
                           lpf_filter_inst_lpf_i_add_271_n1);
   lpf_filter_inst_lpf_i_add_271_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_204_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_133_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_n1, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_2_port, S => 
                           lpf_filter_inst_lpf_i_n67);
   lpf_filter_inst_lpf_i_add_271_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_205_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_134_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_2_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_3_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_2_port);
   lpf_filter_inst_lpf_i_add_271_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_206_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_135_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_3_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_4_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_3_port);
   lpf_filter_inst_lpf_i_add_271_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_207_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_136_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_4_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_5_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_4_port);
   lpf_filter_inst_lpf_i_add_271_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_208_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_137_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_5_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_6_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_5_port);
   lpf_filter_inst_lpf_i_add_271_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_209_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_138_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_6_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_7_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_6_port);
   lpf_filter_inst_lpf_i_add_271_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_210_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_139_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_7_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_8_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_7_port);
   lpf_filter_inst_lpf_i_add_271_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_211_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_140_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_8_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_9_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_8_port);
   lpf_filter_inst_lpf_i_add_271_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_212_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_141_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_9_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_10_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_9_port);
   lpf_filter_inst_lpf_i_add_271_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_213_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_142_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_10_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_11_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_10_port);
   lpf_filter_inst_lpf_i_add_271_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_214_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_143_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_11_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_carry_12_port, S => 
                           lpf_filter_inst_lpf_i_pair11_17_11_port);
   lpf_filter_inst_lpf_i_add_271_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_214_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_143_port, CI => 
                           lpf_filter_inst_lpf_i_add_271_carry_12_port, CO => 
                           lpf_filter_inst_lpf_i_add_271_n_1303, S => 
                           lpf_filter_inst_lpf_i_pair11_17_12_port);
   lpf_filter_inst_lpf_i_add_268_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_84_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_251_port, Z => 
                           lpf_filter_inst_lpf_i_pair7_21_0_port);
   lpf_filter_inst_lpf_i_add_268_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_84_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_251_port, Z => 
                           lpf_filter_inst_lpf_i_add_268_n1);
   lpf_filter_inst_lpf_i_add_268_U1_12 : EXOR3D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_262_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_95_port, A3 => 
                           lpf_filter_inst_lpf_i_add_268_carry_12_port, Z => 
                           lpf_filter_inst_lpf_i_pair7_21_12_port);
   lpf_filter_inst_lpf_i_add_268_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_252_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_85_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_n1, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_2_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_1_port);
   lpf_filter_inst_lpf_i_add_268_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_253_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_86_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_2_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_3_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_2_port);
   lpf_filter_inst_lpf_i_add_268_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_254_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_87_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_3_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_4_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_3_port);
   lpf_filter_inst_lpf_i_add_268_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_255_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_88_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_4_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_5_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_4_port);
   lpf_filter_inst_lpf_i_add_268_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_256_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_89_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_5_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_6_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_5_port);
   lpf_filter_inst_lpf_i_add_268_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_257_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_90_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_6_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_7_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_6_port);
   lpf_filter_inst_lpf_i_add_268_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_258_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_91_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_7_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_8_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_7_port);
   lpf_filter_inst_lpf_i_add_268_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_259_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_92_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_8_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_9_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_8_port);
   lpf_filter_inst_lpf_i_add_268_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_260_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_93_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_9_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_10_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_9_port);
   lpf_filter_inst_lpf_i_add_268_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_261_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_94_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_10_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_11_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_10_port);
   lpf_filter_inst_lpf_i_add_268_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_262_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_95_port, CI => 
                           lpf_filter_inst_lpf_i_add_268_carry_11_port, CO => 
                           lpf_filter_inst_lpf_i_add_268_carry_12_port, S => 
                           lpf_filter_inst_lpf_i_pair7_21_11_port);
   lpf_filter_inst_lpf_i_add_264_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_12_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_323_port, Z => 
                           lpf_filter_inst_lpf_i_pair1_27_0_port);
   lpf_filter_inst_lpf_i_add_264_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_12_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_323_port, Z => 
                           lpf_filter_inst_lpf_i_add_264_n1);
   lpf_filter_inst_lpf_i_add_264_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_324_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_13_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_n1, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_2_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_1_port);
   lpf_filter_inst_lpf_i_add_264_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_325_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_14_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_2_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_3_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_2_port);
   lpf_filter_inst_lpf_i_add_264_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_326_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_15_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_3_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_4_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_3_port);
   lpf_filter_inst_lpf_i_add_264_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_327_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_16_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_4_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_5_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_4_port);
   lpf_filter_inst_lpf_i_add_264_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_328_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_17_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_5_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_6_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_5_port);
   lpf_filter_inst_lpf_i_add_264_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_329_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_18_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_6_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_7_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_6_port);
   lpf_filter_inst_lpf_i_add_264_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_330_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_19_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_7_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_8_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_7_port);
   lpf_filter_inst_lpf_i_add_264_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_331_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_20_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_8_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_9_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_8_port);
   lpf_filter_inst_lpf_i_add_264_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_332_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_21_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_9_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_10_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_9_port);
   lpf_filter_inst_lpf_i_add_264_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_333_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_22_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_10_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_11_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_10_port);
   lpf_filter_inst_lpf_i_add_264_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_334_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_23_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_11_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_carry_12_port, S => 
                           lpf_filter_inst_lpf_i_pair1_27_11_port);
   lpf_filter_inst_lpf_i_add_264_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_334_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_23_port, CI => 
                           lpf_filter_inst_lpf_i_add_264_carry_12_port, CO => 
                           lpf_filter_inst_lpf_i_add_264_n_1298, S => 
                           lpf_filter_inst_lpf_i_pair1_27_12_port);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_0_port, A2 => 
                           mixer_out_i_0_port, Z => 
                           lpf_filter_inst_lpf_i_pair0_28_0);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_0_port, A2 => 
                           mixer_out_i_0_port, Z => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_n1);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_12 : EXOR3D1 port map( A1 => 
                           mixer_out_i_11_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_11_port, A3 => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_12_port, Z 
                           => lpf_filter_inst_lpf_i_pair0_28_12);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_1 : ADFULD1 port map( A => 
                           mixer_out_i_1_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_1_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_2_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_1);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_2 : ADFULD1 port map( A => 
                           mixer_out_i_2_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_2_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_2);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_3 : ADFULD1 port map( A => 
                           mixer_out_i_3_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_3_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_3);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_4 : ADFULD1 port map( A => 
                           mixer_out_i_4_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_4_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_4);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_5 : ADFULD1 port map( A => 
                           mixer_out_i_5_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_5_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_5);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_6 : ADFULD1 port map( A => 
                           mixer_out_i_6_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_6_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_6);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_7 : ADFULD1 port map( A => 
                           mixer_out_i_7_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_7_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_7);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_8 : ADFULD1 port map( A => 
                           mixer_out_i_8_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_8_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_8);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_9 : ADFULD1 port map( A => 
                           mixer_out_i_9_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_9_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_9);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_10 : ADFULD1 port map( A => 
                           mixer_out_i_10_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_10_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_10);
   lpf_filter_inst_lpf_i_add_5_root_add_292_U1_11 : ADFULD1 port map( A => 
                           mixer_out_i_11_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_11_port, CI => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_5_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_pair0_28_11);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair12_16_1_port, A2 => 
                           lpf_filter_inst_lpf_i_pair1_27_0_port, Z => 
                           lpf_filter_inst_lpf_i_t0_1_1);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair12_16_1_port, A2 => 
                           lpf_filter_inst_lpf_i_pair1_27_0_port, Z => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_n1);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_14 : EXOR3D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair1_27_12_port, A2 => 
                           lpf_filter_inst_lpf_i_n1, A3 => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_14_port, Z 
                           => lpf_filter_inst_lpf_i_t0_1_14);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_1_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_2_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_2);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_2_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_3_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_3);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_3_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_4_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_4);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_4_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_5_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_5);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_5_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_6_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_6);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_6_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_7_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_7);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_7_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_8_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_8);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_8_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_9_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_9);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_9_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_10_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_10);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_10_port, B => 
                           lpf_filter_inst_lpf_i_pair12_16_11_port, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_11);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_11_port, B => 
                           lpf_filter_inst_lpf_i_n1, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_12);
   lpf_filter_inst_lpf_i_add_4_root_add_292_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair1_27_12_port, B => 
                           lpf_filter_inst_lpf_i_n1, CI => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_4_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_t0_1_13);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_p141_1_2_port, A2 => 
                           lpf_filter_inst_lpf_i_t11_14_0_port, Z => 
                           lpf_filter_inst_lpf_i_n156);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_p141_1_2_port, A2 => 
                           lpf_filter_inst_lpf_i_t11_14_0_port, Z => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_n1);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_1_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_3_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_n155);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_2_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_4_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_n154);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_3_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_5_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_n153);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_4_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_6_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_n152);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_5_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_7_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_n151);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_6_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_8_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_n150);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_7_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_9_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_n149);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_8_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_10_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_n148);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_9_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_11_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_n147);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_10_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_12_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_n146);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_11_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_13_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_n145);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_12_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_14_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_n144);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_13_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_15_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_n143);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_14_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_16_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_n142);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_15_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_17_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_i_n141);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_16_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_19_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_i_n140);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_20 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_17_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_19_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_i_n139);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_21 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_18_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_19_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_i_n138);
   lpf_filter_inst_lpf_i_add_7_root_add_292_U1_22 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_18_port, B => 
                           lpf_filter_inst_lpf_i_p141_1_19_port, CI => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_7_root_add_292_n_1017, S 
                           => lpf_filter_inst_lpf_i_n137);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_3_port, A2 => 
                           lpf_filter_inst_lpf_i_t3_7_1_port, Z => 
                           lpf_filter_inst_lpf_i_n135);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_3_port, A2 => 
                           lpf_filter_inst_lpf_i_t3_7_1_port, Z => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_n1);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_2_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_4_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_n134);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_3_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_5_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_n133);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_4_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_6_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_n132);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_5_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_7_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_n131);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_6_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_8_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_n130);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_7_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_9_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_n129);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_8_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_10_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_n128);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_9_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_11_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_n127);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_10_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_12_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_n126);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_11_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_13_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_n125);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_12_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_14_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_n124);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_13_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_15_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_n123);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_14_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_16_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_n122);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_15_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_17_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_n121);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_15_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_18_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_i_n120);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_15_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_19_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_i_n119);
   lpf_filter_inst_lpf_i_add_8_root_add_292_U1_20 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t3_7_15_port, B => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_19_port, CI => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_8_root_add_292_n_1027, S 
                           => lpf_filter_inst_lpf_i_n118);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_p206_3_3_port, A2 => 
                           lpf_filter_inst_lpf_i_n117, Z => 
                           lpf_filter_inst_lpf_i_t12_13_4);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_p206_3_3_port, A2 => 
                           lpf_filter_inst_lpf_i_n117, Z => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_n1);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_1_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_4_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_5);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_2_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_5_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_6);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_3_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_6_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_7);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_4_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_7_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_8);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_5_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_8_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_9);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_6_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_9_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_10);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_7_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_10_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_11);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_8_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_11_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_12);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_9_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_12_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_13);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_10_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_13_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_14);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair12_16_11_port, B => 
                           lpf_filter_inst_lpf_i_p206_3_14_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_15);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n1, B => 
                           lpf_filter_inst_lpf_i_p206_3_15_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_16);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n1, B => 
                           lpf_filter_inst_lpf_i_p206_3_16_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_17);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n1, B => 
                           lpf_filter_inst_lpf_i_p206_3_17_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_18);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n1, B => 
                           lpf_filter_inst_lpf_i_p206_3_18_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_19);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_20 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n1, B => 
                           lpf_filter_inst_lpf_i_p206_3_19_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_20);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_21 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n1, B => 
                           lpf_filter_inst_lpf_i_p206_3_20_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_i_t12_13_21);
   lpf_filter_inst_lpf_i_add_6_root_add_292_U1_22 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n1, B => 
                           lpf_filter_inst_lpf_i_p206_3_20_port, CI => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_6_root_add_292_n_1036, S 
                           => lpf_filter_inst_lpf_i_t12_13_22);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U2 : EXOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_i_n117, A2 => 
                           lpf_filter_inst_lpf_i_p206_1_3, Z => 
                           lpf_filter_inst_lpf_i_n181);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1 : AND2D1 port map( A1
                           => lpf_filter_inst_lpf_i_n117, A2 => 
                           lpf_filter_inst_lpf_i_p206_1_3, Z => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_n1);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_2 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_t12_13_2, B => 
                           lpf_filter_inst_lpf_i_n157, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_n1, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_n180);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_3 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_t12_13_3, B => 
                           lpf_filter_inst_lpf_i_n156, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_n179);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_4 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_t12_13_4, B => 
                           lpf_filter_inst_lpf_i_n155, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_n178);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_5 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_t12_13_5, B => 
                           lpf_filter_inst_lpf_i_n154, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_n177);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_6 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_t12_13_6, B => 
                           lpf_filter_inst_lpf_i_n153, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_n176);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_7 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_t12_13_7, B => 
                           lpf_filter_inst_lpf_i_n152, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_n175);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_8 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_t12_13_8, B => 
                           lpf_filter_inst_lpf_i_n151, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_n174);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_9 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_t12_13_9, B => 
                           lpf_filter_inst_lpf_i_n150, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_n173);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_10 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_10, B => 
                           lpf_filter_inst_lpf_i_n149, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_n172);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_11 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_11, B => 
                           lpf_filter_inst_lpf_i_n148, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_n171);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_12 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_12, B => 
                           lpf_filter_inst_lpf_i_n147, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_n170);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_13 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_13, B => 
                           lpf_filter_inst_lpf_i_n146, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_n169);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_14 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_14, B => 
                           lpf_filter_inst_lpf_i_n145, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_n168);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_15 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_15, B => 
                           lpf_filter_inst_lpf_i_n144, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_n167);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_16 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_16, B => 
                           lpf_filter_inst_lpf_i_n143, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_n166);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_17 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_17, B => 
                           lpf_filter_inst_lpf_i_n142, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_n165);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_18 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_18, B => 
                           lpf_filter_inst_lpf_i_n141, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_i_n164);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_19 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_19, B => 
                           lpf_filter_inst_lpf_i_n140, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_i_n163);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_20 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_20, B => 
                           lpf_filter_inst_lpf_i_n139, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_i_n162);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_21 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_21, B => 
                           lpf_filter_inst_lpf_i_n138, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_i_n161);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_22 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_22, B => 
                           lpf_filter_inst_lpf_i_n137, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_23_port, S 
                           => lpf_filter_inst_lpf_i_n160);
   lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_U1_23 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_t12_13_22, B => 
                           lpf_filter_inst_lpf_i_n137, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_carry_23_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_0_root_add_292_n_1042, S 
                           => lpf_filter_inst_lpf_i_n159);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U17 : EXOR2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n15, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n16, Z 
                           => lpf_filter_inst_lpf_i_n92);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U16 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_2, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n14);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U15 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_1, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n15);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U14 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_3, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n13);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U13 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_n117, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n16);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U12 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_14, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U11 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_13, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n3);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U10 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_12, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n4);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U9 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_11, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n5);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U8 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_10, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n6);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U7 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_9, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n7);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U6 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_8, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n8);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U5 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_7, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n9);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U4 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_6, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n10);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U3 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_5, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n11);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_t0_1_4, Z => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n12);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U1 : AND2D1 port map( A1
                           => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n15, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n16, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n1);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_2 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n136, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n14, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n1, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_n91);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_3 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n135, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n13, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_n90);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_4 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n134, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n12, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_n89);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_5 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n133, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n11, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_n88);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_6 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n132, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n10, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_n87);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_7 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n131, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n9, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_n86);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_8 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n130, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n8, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_n85);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_9 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n129, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n7, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_n84);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_10 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n128, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n6, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_n83);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_11 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n127, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n5, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_n194);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_12 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n126, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n4, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_n193);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_13 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n125, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n3, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_n192);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_14 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n124, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_n191);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_15 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n123, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_n190);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_16 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n122, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_n189);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_17 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n121, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_n188);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_18 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n120, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_i_n187);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_19 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n119, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_i_n186);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_20 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n118, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_i_n185);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_21 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n118, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_i_n184);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_22 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n118, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_23_port, S 
                           => lpf_filter_inst_lpf_i_n183);
   lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_U2_23 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n118, B => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_carry_23_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_3_root_sub_0_root_add_292_n_1047, S 
                           => lpf_filter_inst_lpf_i_n182);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U2 : EXOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_i_n181, A2 => 
                           lpf_filter_inst_lpf_i_n92, Z => 
                           lpf_filter_inst_lpf_i_n116);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1 : AND2D1 port map( A1
                           => lpf_filter_inst_lpf_i_n181, A2 => 
                           lpf_filter_inst_lpf_i_n92, Z => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_n1);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_2 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n91, B => 
                           lpf_filter_inst_lpf_i_n180, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_n1, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_n115);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_3 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n90, B => 
                           lpf_filter_inst_lpf_i_n179, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_n114);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_4 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n89, B => 
                           lpf_filter_inst_lpf_i_n178, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_n113);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_5 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n88, B => 
                           lpf_filter_inst_lpf_i_n177, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_n112);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_6 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n87, B => 
                           lpf_filter_inst_lpf_i_n176, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_n111);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_7 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n86, B => 
                           lpf_filter_inst_lpf_i_n175, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_n110);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_8 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n85, B => 
                           lpf_filter_inst_lpf_i_n174, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_n109);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_9 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_i_n84, B => 
                           lpf_filter_inst_lpf_i_n173, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_n108);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_10 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n83, B => 
                           lpf_filter_inst_lpf_i_n172, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_n107);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_11 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n194, B => 
                           lpf_filter_inst_lpf_i_n171, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_n106);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_12 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n193, B => 
                           lpf_filter_inst_lpf_i_n170, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_n105);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_13 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n192, B => 
                           lpf_filter_inst_lpf_i_n169, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_n104);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_14 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n191, B => 
                           lpf_filter_inst_lpf_i_n168, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_n103);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_15 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n190, B => 
                           lpf_filter_inst_lpf_i_n167, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_n102);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_16 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n189, B => 
                           lpf_filter_inst_lpf_i_n166, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_n101);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_17 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n188, B => 
                           lpf_filter_inst_lpf_i_n165, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_n100);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_18 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n187, B => 
                           lpf_filter_inst_lpf_i_n164, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_i_n99);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_19 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n186, B => 
                           lpf_filter_inst_lpf_i_n163, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_i_n98);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_20 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n185, B => 
                           lpf_filter_inst_lpf_i_n162, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_i_n97);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_21 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n184, B => 
                           lpf_filter_inst_lpf_i_n161, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_i_n96);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_22 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n183, B => 
                           lpf_filter_inst_lpf_i_n160, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_23_port, S 
                           => lpf_filter_inst_lpf_i_n95);
   lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_U1_23 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n182, B => 
                           lpf_filter_inst_lpf_i_n159, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_carry_23_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_0_root_add_292_n_1051, S 
                           => lpf_filter_inst_lpf_i_n94);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U30 : NOR2M1D1 port map(
                           A1 => lpf_filter_inst_lpf_i_pair0_28_0, A2 => 
                           lpf_filter_inst_lpf_i_n117, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n28);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U29 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n28, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n7, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n29);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U28 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n28, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n7, 
                           B1 => lpf_filter_inst_lpf_i_pair0_28_1, B2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n29, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n26);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U27 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_i_n115, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n26, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n27);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U26 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n26, 
                           B2 => lpf_filter_inst_lpf_i_n115, A1 => 
                           lpf_filter_inst_lpf_i_pair0_28_2, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n27, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n24);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U25 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n24, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n6, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n25);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U24 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n24, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n6, 
                           B1 => lpf_filter_inst_lpf_i_pair0_28_3, B2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n25, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n22);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U23 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_i_n113, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n22, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n23);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U22 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n22, 
                           B2 => lpf_filter_inst_lpf_i_n113, A1 => 
                           lpf_filter_inst_lpf_i_pair0_28_4, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n23, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n20);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U21 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n20, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n5, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n21);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U20 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n20, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n5, 
                           B1 => lpf_filter_inst_lpf_i_pair0_28_5, B2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n21, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n18);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U19 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_i_n111, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n18, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n19);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U18 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n18, 
                           B2 => lpf_filter_inst_lpf_i_n111, A1 => 
                           lpf_filter_inst_lpf_i_pair0_28_6, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n19, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n16);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U17 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n16, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n4, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n17);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U16 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n16, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n4, 
                           B1 => lpf_filter_inst_lpf_i_pair0_28_7, B2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n17, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n14);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U15 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_i_n109, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n14, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n15);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U14 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n14, 
                           B2 => lpf_filter_inst_lpf_i_n109, A1 => 
                           lpf_filter_inst_lpf_i_pair0_28_8, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n15, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n12);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U13 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n12, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n3, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n13);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U12 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n12, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n3, 
                           B1 => lpf_filter_inst_lpf_i_pair0_28_9, B2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n13, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n10);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U11 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_i_n107, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n10, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n11);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U10 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n10, 
                           B2 => lpf_filter_inst_lpf_i_n107, A1 => 
                           lpf_filter_inst_lpf_i_pair0_28_10, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n11, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n8);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U9 : AND2D1 port map( A1
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n8, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n2, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n9);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U8 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n8, 
                           A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n2, 
                           B1 => lpf_filter_inst_lpf_i_pair0_28_11, B2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n9, Z 
                           => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_12_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U7 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_pair0_28_12, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U6 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_n108, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n3);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U5 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_n110, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n4);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U4 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_n112, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n5);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U3 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_n114, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n6);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_n116, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n7);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U1 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_i_n106, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n2);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_12 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n105, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_13_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_12_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_13 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n104, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_14_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_13_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_14 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n103, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_15_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_14_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_15 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n102, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_16_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_15_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_16 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n101, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_17_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_16_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_17 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n100, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_18_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_17_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_18 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n99, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_19_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_18_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_19 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n98, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_20_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_19_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_20 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n97, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_21_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_20_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_21 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n96, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_22_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_21_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_22 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n95, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_23_port, S 
                           => 
                           lpf_filter_inst_lpf_i_t0_1_3_4_5_7_8_9_11_12_13_14_22_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_U2_23 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_i_n94, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_carry_23_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_0_root_add_292_n_1066, S 
                           => filter_out_i_4_port);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_p206_2_3_port, A2 => 
                           lpf_filter_inst_lpf_i_p206_1_3, Z => 
                           lpf_filter_inst_lpf_i_p206_1_6);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_p206_2_3_port, A2 => 
                           lpf_filter_inst_lpf_i_p206_1_3, Z => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_n1);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_1_4, B => 
                           lpf_filter_inst_lpf_i_p206_2_4_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_n1, CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_7);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_2_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_5_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_8);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_3_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_6_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_9);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_4_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_7_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_10);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_5_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_8_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_11);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_6_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_9_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_12);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_7_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_10_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_13);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_8_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_11_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_14);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_9_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_12_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_15);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_10_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_13_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_16);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair13_15_11_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_14_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_17);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_2_15_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_15_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_19_port, S 
                           => lpf_filter_inst_lpf_i_p206_1_18);
   lpf_filter_inst_lpf_i_add_1_root_add_285_U1_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_p206_2_15_port, B => 
                           lpf_filter_inst_lpf_i_p206_2_15_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_285_n_1143, S 
                           => lpf_filter_inst_lpf_i_p206_1_19);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_60_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_275_port, Z => 
                           lpf_filter_inst_lpf_i_pair4_24_0);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_60_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_275_port, Z => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_n1);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_276_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_61_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_n1, CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_2_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_1);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_277_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_62_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_2);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_278_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_63_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_3);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_279_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_64_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_4);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_280_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_65_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_5);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_281_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_66_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_6);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_282_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_67_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_7);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_283_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_68_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_8);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_284_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_69_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_9);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_285_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_70_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_10);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_286_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_71_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_pair4_24_11);
   lpf_filter_inst_lpf_i_add_2_root_sub_287_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_286_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_71_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_sub_287_n_1254, S 
                           => lpf_filter_inst_lpf_i_pair4_24_12);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_48_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_287_port, Z => 
                           lpf_filter_inst_lpf_i_pair5_23_0);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_48_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_287_port, Z => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_n1);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_288_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_49_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_n1, CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_2_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_1);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_289_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_50_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_2);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_290_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_51_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_3);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_291_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_52_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_4);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_292_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_53_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_5);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_293_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_54_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_6);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_294_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_55_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_7);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_295_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_56_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_8);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_296_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_57_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_9);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_297_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_58_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_10);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_298_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_59_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_pair5_23_11);
   lpf_filter_inst_lpf_i_add_3_root_sub_287_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_298_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_59_port, CI => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_3_root_sub_287_n_1257, S 
                           => lpf_filter_inst_lpf_i_pair5_23_12);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair4_24_0, A2 => 
                           lpf_filter_inst_lpf_i_pair5_23_0, Z => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_3_port);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair4_24_0, A2 => 
                           lpf_filter_inst_lpf_i_pair5_23_0, Z => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_n1);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_1, B => 
                           lpf_filter_inst_lpf_i_pair4_24_1, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_n1, CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_2_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_4_port);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_2, B => 
                           lpf_filter_inst_lpf_i_pair4_24_2, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_2);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_3, B => 
                           lpf_filter_inst_lpf_i_pair4_24_3, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_3);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_4, B => 
                           lpf_filter_inst_lpf_i_pair4_24_4, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_4);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_5, B => 
                           lpf_filter_inst_lpf_i_pair4_24_5, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_5);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_6, B => 
                           lpf_filter_inst_lpf_i_pair4_24_6, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_6);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_7, B => 
                           lpf_filter_inst_lpf_i_pair4_24_7, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_7);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_8, B => 
                           lpf_filter_inst_lpf_i_pair4_24_8, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_9, B => 
                           lpf_filter_inst_lpf_i_pair4_24_9, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_9);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_10, B => 
                           lpf_filter_inst_lpf_i_pair4_24_10, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_10);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_11, B => 
                           lpf_filter_inst_lpf_i_pair4_24_11, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_11);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_12, B => 
                           lpf_filter_inst_lpf_i_pair4_24_12, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_12);
   lpf_filter_inst_lpf_i_add_1_root_sub_287_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair5_23_12, B => 
                           lpf_filter_inst_lpf_i_pair4_24_12, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_287_n_1260, S 
                           => lpf_filter_inst_lpf_i_t4_5_13);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U17 : EXNOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n15, A2 => 
                           lpf_filter_inst_lpf_i_t4_5_2, Z => 
                           lpf_filter_inst_lpf_i_t4_5_8_9_5_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U16 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_0_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n15);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U15 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_13_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n2);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U14 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_2, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n1);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U13 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_10_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n5);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U12 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_9_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n6);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U11 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_8_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n7);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U10 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_7_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n8);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U9 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_6_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n9);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U8 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_5_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n10);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U7 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_4_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n11);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U6 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_3_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n12);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U5 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_2_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n13);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U4 : NAN2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t8_9_0_port, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n1, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_3_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U3 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_1_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n14);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_12_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n3);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U1 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t8_9_11_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n4);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_3, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n14, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_6_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_4, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n13, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_7_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_5, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n12, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_8_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_6, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n11, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_9_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_7, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n10, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_10_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_8, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n9, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_11_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_9, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n8, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_12_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_10, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n7, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_13_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_11, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n6, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_14_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_12, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n5, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_15_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_13, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n4, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_16_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_13, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n3, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_17_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_13, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n2, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_18_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_287_U2_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_t4_5_13, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n2, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_287_n_1265, S 
                           => lpf_filter_inst_lpf_i_t4_5_8_9_19_port);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t11_14_0_port, A2 => 
                           lpf_filter_inst_lpf_i_pair11_17_2_port, Z => 
                           lpf_filter_inst_lpf_i_n66);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_t11_14_0_port, A2 => 
                           lpf_filter_inst_lpf_i_pair11_17_2_port, Z => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_n1);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_3_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_168_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_n1, CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_n65);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_4_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_169_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_n64);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_5_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_170_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_n63);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_6_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_171_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_n82);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_7_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_172_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_n81);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_8_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_173_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_n80);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_9_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_174_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_n79);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_10_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_175_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_n78);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_11_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_176_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_n77);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_12_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_177_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_n76);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_12_port, B => 
                           lpf_filter_inst_lpf_i_p232_2_17, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_n75);
   lpf_filter_inst_lpf_i_add_2_root_add_286_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair11_17_12_port, B => 
                           lpf_filter_inst_lpf_i_p232_2_17, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_286_n_1180, S 
                           => lpf_filter_inst_lpf_i_n62);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U22 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n19, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n20, Z => 
                           lpf_filter_inst_lpf_i_t11_14_1_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U21 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n18, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n2, Z => 
                           lpf_filter_inst_lpf_i_t11_14_2_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U20 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_1, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n19);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U19 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_t11_14_0_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n20);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U18 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_5, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n15);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U17 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_3, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n17);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U16 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n19, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n20, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n2);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U15 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_2, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n18);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U14 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_17, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n3);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U13 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_17, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n4);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U12 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_17, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n5);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U11 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_17, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n6);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U10 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_17, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n7);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U9 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_12, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n8);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U8 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_11, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n9);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U7 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_10, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n10);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U6 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_9, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n11);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U5 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_8, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n12);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U4 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_7, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n13);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U3 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_6, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n14);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_p232_2_4, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n16);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n18, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n2, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n1);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n74, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n17, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n1, CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_3_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n67, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n16, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_4_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n66, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n15, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_5_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n65, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n14, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_6_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n64, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n13, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_7_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n63, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n12, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_8_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n82, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n11, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_9_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n81, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n10, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_10_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n80, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n9, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_11_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n79, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n8, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_12_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n78, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n7, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_13_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n77, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n6, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_14_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n76, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n5, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_16_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_15_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n75, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n4, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_17_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_16_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n62, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n3, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_18_port, S 
                           => lpf_filter_inst_lpf_i_t11_14_17_port);
   lpf_filter_inst_lpf_i_sub_0_root_add_286_U2_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_n62, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n3, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_add_286_n_1186, S 
                           => lpf_filter_inst_lpf_i_t11_14_18_port);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_108_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_227_port, Z => 
                           lpf_filter_inst_lpf_i_pair8_20_0);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_108_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_227_port, Z => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_n1);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_228_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_109_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_n1, CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_2_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_1);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_229_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_110_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_2);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_230_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_111_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_3);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_231_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_112_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_4);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_232_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_113_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_5);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_233_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_114_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_6);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_234_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_115_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_7);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_235_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_116_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_8);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_236_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_117_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_9);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_237_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_118_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_10);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_238_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_119_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_pair8_20_11);
   lpf_filter_inst_lpf_i_add_1_root_add_277_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_238_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_119_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_add_277_n_1282, S 
                           => lpf_filter_inst_lpf_i_pair8_20_12);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_96_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_239_port, Z => 
                           lpf_filter_inst_lpf_i_pair9_19_0);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_96_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_239_port, Z => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_n1);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_240_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_97_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_n1, CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_2_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_1);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_241_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_98_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_2);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_242_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_99_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_3);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_243_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_100_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_4);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_244_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_101_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_5);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_245_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_102_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_6);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_246_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_103_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_7);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_247_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_104_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_8);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_248_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_105_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_9);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_249_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_106_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_10);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_250_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_107_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_pair9_19_11);
   lpf_filter_inst_lpf_i_add_2_root_add_277_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_250_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_107_port, CI => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_2_root_add_277_n_1285, S 
                           => lpf_filter_inst_lpf_i_pair9_19_12);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair8_20_0, A2 => 
                           lpf_filter_inst_lpf_i_pair9_19_0, Z => 
                           lpf_filter_inst_lpf_i_t8_9_0_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair8_20_0, A2 => 
                           lpf_filter_inst_lpf_i_pair9_19_0, Z => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_n1);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_13 : EXOR3D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair9_19_12, A2 => 
                           lpf_filter_inst_lpf_i_pair8_20_12, A3 => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_13_port, Z 
                           => lpf_filter_inst_lpf_i_t8_9_13_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_1, B => 
                           lpf_filter_inst_lpf_i_pair8_20_1, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_n1, CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_2_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_1_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_2, B => 
                           lpf_filter_inst_lpf_i_pair8_20_2, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_2_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_3, B => 
                           lpf_filter_inst_lpf_i_pair8_20_3, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_3_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_4, B => 
                           lpf_filter_inst_lpf_i_pair8_20_4, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_4_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_5, B => 
                           lpf_filter_inst_lpf_i_pair8_20_5, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_5_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_6, B => 
                           lpf_filter_inst_lpf_i_pair8_20_6, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_6_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_7, B => 
                           lpf_filter_inst_lpf_i_pair8_20_7, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_7_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_8, B => 
                           lpf_filter_inst_lpf_i_pair8_20_8, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_8_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_9, B => 
                           lpf_filter_inst_lpf_i_pair8_20_9, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_9_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_10, B => 
                           lpf_filter_inst_lpf_i_pair8_20_10, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_10_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_11, B => 
                           lpf_filter_inst_lpf_i_pair8_20_11, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_11_port);
   lpf_filter_inst_lpf_i_add_0_root_add_277_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair9_19_12, B => 
                           lpf_filter_inst_lpf_i_pair8_20_12, CI => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_0_root_add_277_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_t8_9_12_port);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_36_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_299_port, Z => 
                           lpf_filter_inst_lpf_i_n136);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_36_port, A2 => 
                           lpf_filter_inst_lpf_i_arx_input_reg_299_port, Z => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_n1);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_300_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_37_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_n1, CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_2_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_1_port);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_301_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_38_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_3_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_2);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_302_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_39_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_3);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_303_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_40_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_4);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_304_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_41_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_5);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_305_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_42_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_6);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_306_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_43_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_7);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_307_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_44_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_8);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_308_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_45_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_9);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_309_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_46_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_10);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_310_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_47_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_pair3_25_11);
   lpf_filter_inst_lpf_i_add_1_root_sub_279_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_arx_input_reg_310_port, B => 
                           lpf_filter_inst_lpf_i_arx_input_reg_47_port, CI => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_add_1_root_sub_279_n_1161, S 
                           => lpf_filter_inst_lpf_i_pair3_25_12);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U16 : EXNOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n14, A2 => 
                           lpf_filter_inst_lpf_i_pair3_25_2, Z => 
                           lpf_filter_inst_lpf_i_t3_7_2_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U15 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_0_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n14);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U14 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_12_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n2);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U13 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_2, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n1);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U12 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_9_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n5);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U11 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_8_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n6);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U10 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_7_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n7);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U9 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_6_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n8);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U8 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_5_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n9);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U7 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_4_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n10);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U6 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_3_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n11);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U5 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_2_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n12);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U4 : NAN2D1 port map( A1 => 
                           lpf_filter_inst_lpf_i_pair7_21_0_port, A2 => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n1, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_3_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U3 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_1_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n13);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_11_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n3);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U1 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair7_21_10_port, Z => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n4);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_3, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n13, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_4_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_3_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_4, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n12, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_5_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_4_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_5, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n11, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_6_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_5_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_6, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n10, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_7_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_6_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_7, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n9, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_8_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_7_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_8, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n8, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_9_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_8_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_9, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n7, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_10_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_9_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_10, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n6, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_11_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_10_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_11, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n5, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_12_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_11_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_12, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n4, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_13_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_12_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_12, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n3, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_14_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_13_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_12, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n2, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_15_port, S 
                           => lpf_filter_inst_lpf_i_t3_7_14_port);
   lpf_filter_inst_lpf_i_sub_0_root_sub_279_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_i_pair3_25_12, B => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n2, CI => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_i_sub_0_root_sub_279_n_1166, S 
                           => lpf_filter_inst_lpf_i_t3_7_15_port);
   lpf_filter_inst_lpf_q_U94 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair13_15_2_port, A2 => 
                           lpf_filter_inst_lpf_q_p206_1_3, Z => 
                           lpf_filter_inst_lpf_q_p206_1_5);
   lpf_filter_inst_lpf_q_U93 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair13_15_2_port, A2 => 
                           lpf_filter_inst_lpf_q_p206_1_3, Z => 
                           lpf_filter_inst_lpf_q_add_284_carry_3);
   lpf_filter_inst_lpf_q_U92 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_n37, A2 => 
                           lpf_filter_inst_lpf_q_n36, Z => 
                           lpf_filter_inst_lpf_q_t12_13_2);
   lpf_filter_inst_lpf_q_U91 : AND2D1 port map( A1 => lpf_filter_inst_lpf_q_n36
                           , A2 => lpf_filter_inst_lpf_q_n37, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_2_port);
   lpf_filter_inst_lpf_q_U90 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_n38, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_2_port, Z 
                           => lpf_filter_inst_lpf_q_t12_13_3);
   lpf_filter_inst_lpf_q_U89 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_2_port, 
                           A2 => lpf_filter_inst_lpf_q_n38, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_3_port);
   lpf_filter_inst_lpf_q_U88 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t11_14_0_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_168_port, Z => 
                           lpf_filter_inst_lpf_q_p232_2_1);
   lpf_filter_inst_lpf_q_U87 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t11_14_0_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_168_port, Z => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_2);
   lpf_filter_inst_lpf_q_U86 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_n50, A2 => 
                           lpf_filter_inst_lpf_q_n49, Z => 
                           lpf_filter_inst_lpf_q_n157);
   lpf_filter_inst_lpf_q_U85 : AND2D1 port map( A1 => lpf_filter_inst_lpf_q_n49
                           , A2 => lpf_filter_inst_lpf_q_n50, Z => 
                           lpf_filter_inst_lpf_q_sub_280_carry_2_port);
   lpf_filter_inst_lpf_q_U84 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_n51, A2 => 
                           lpf_filter_inst_lpf_q_sub_280_carry_2_port, Z => 
                           lpf_filter_inst_lpf_q_p141_1_2_port);
   lpf_filter_inst_lpf_q_U83 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_280_carry_2_port, A2 => 
                           lpf_filter_inst_lpf_q_n51, Z => 
                           lpf_filter_inst_lpf_q_sub_280_carry_3_port);
   lpf_filter_inst_lpf_q_U82 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_n52, A2 => 
                           lpf_filter_inst_lpf_q_sub_280_carry_3_port, Z => 
                           lpf_filter_inst_lpf_q_p141_1_3_port);
   lpf_filter_inst_lpf_q_U81 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_280_carry_3_port, A2 => 
                           lpf_filter_inst_lpf_q_n52, Z => 
                           lpf_filter_inst_lpf_q_sub_280_carry_4_port);
   lpf_filter_inst_lpf_q_U80 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_n53, A2 => 
                           lpf_filter_inst_lpf_q_sub_280_carry_4_port, Z => 
                           lpf_filter_inst_lpf_q_p141_1_4_port);
   lpf_filter_inst_lpf_q_U79 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_280_carry_4_port, A2 => 
                           lpf_filter_inst_lpf_q_n53, Z => 
                           lpf_filter_inst_lpf_q_sub_280_carry_5_port);
   lpf_filter_inst_lpf_q_U78 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_n54, A2 => 
                           lpf_filter_inst_lpf_q_sub_280_carry_5_port, Z => 
                           lpf_filter_inst_lpf_q_p141_1_5_port);
   lpf_filter_inst_lpf_q_U77 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_280_carry_5_port, A2 => 
                           lpf_filter_inst_lpf_q_n54, Z => 
                           lpf_filter_inst_lpf_q_sub_280_carry_6_port);
   lpf_filter_inst_lpf_q_U76 : TIELO port map( Z => 
                           lpf_filter_inst_lpf_q_net5308);
   lpf_filter_inst_lpf_q_U75 : INVD1 port map( A => rstn, Z => 
                           lpf_filter_inst_lpf_q_n3);
   lpf_filter_inst_lpf_q_U74 : BUFD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_12_port, Z => 
                           lpf_filter_inst_lpf_q_n1);
   lpf_filter_inst_lpf_q_U73 : BUFD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_178_port, Z => 
                           lpf_filter_inst_lpf_q_p232_2_17);
   lpf_filter_inst_lpf_q_U72 : INVD1 port map( A => lpf_filter_inst_lpf_q_n3, Z
                           => lpf_filter_inst_lpf_q_n2);
   lpf_filter_inst_lpf_q_U71 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_2_port, Z => 
                           lpf_filter_inst_lpf_q_n38);
   lpf_filter_inst_lpf_q_U70 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_3, Z => 
                           lpf_filter_inst_lpf_q_n36);
   lpf_filter_inst_lpf_q_U69 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_5_port, Z => 
                           lpf_filter_inst_lpf_q_n54);
   lpf_filter_inst_lpf_q_U68 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_4_port, Z => 
                           lpf_filter_inst_lpf_q_n53);
   lpf_filter_inst_lpf_q_U67 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_3_port, Z => 
                           lpf_filter_inst_lpf_q_n52);
   lpf_filter_inst_lpf_q_U66 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_2_port, Z => 
                           lpf_filter_inst_lpf_q_n51);
   lpf_filter_inst_lpf_q_U65 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_4, Z => 
                           lpf_filter_inst_lpf_q_n37);
   lpf_filter_inst_lpf_q_U64 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_1_port, Z => 
                           lpf_filter_inst_lpf_q_n50);
   lpf_filter_inst_lpf_q_U63 : INVD1 port map( A => lpf_filter_inst_lpf_q_n117,
                           Z => lpf_filter_inst_lpf_q_n49);
   lpf_filter_inst_lpf_q_U62 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_11_port, Z => 
                           lpf_filter_inst_lpf_q_n47);
   lpf_filter_inst_lpf_q_U61 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_10_port, Z => 
                           lpf_filter_inst_lpf_q_n46);
   lpf_filter_inst_lpf_q_U60 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_9_port, Z => 
                           lpf_filter_inst_lpf_q_n45);
   lpf_filter_inst_lpf_q_U59 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_8_port, Z => 
                           lpf_filter_inst_lpf_q_n44);
   lpf_filter_inst_lpf_q_U58 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_7_port, Z => 
                           lpf_filter_inst_lpf_q_n43);
   lpf_filter_inst_lpf_q_U57 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_6_port, Z => 
                           lpf_filter_inst_lpf_q_n42);
   lpf_filter_inst_lpf_q_U56 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_5_port, Z => 
                           lpf_filter_inst_lpf_q_n41);
   lpf_filter_inst_lpf_q_U55 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_11_port, Z => 
                           lpf_filter_inst_lpf_q_n60);
   lpf_filter_inst_lpf_q_U54 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_10_port, Z => 
                           lpf_filter_inst_lpf_q_n59);
   lpf_filter_inst_lpf_q_U53 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_9_port, Z => 
                           lpf_filter_inst_lpf_q_n58);
   lpf_filter_inst_lpf_q_U52 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_8_port, Z => 
                           lpf_filter_inst_lpf_q_n57);
   lpf_filter_inst_lpf_q_U51 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_4_port, Z => 
                           lpf_filter_inst_lpf_q_n40);
   lpf_filter_inst_lpf_q_U50 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_7_port, Z => 
                           lpf_filter_inst_lpf_q_n56);
   lpf_filter_inst_lpf_q_U49 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_3_port, Z => 
                           lpf_filter_inst_lpf_q_n39);
   lpf_filter_inst_lpf_q_U48 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_6_port, Z => 
                           lpf_filter_inst_lpf_q_n55);
   lpf_filter_inst_lpf_q_U47 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_2_15_port, Z => 
                           lpf_filter_inst_lpf_q_n48);
   lpf_filter_inst_lpf_q_U46 : INVD1 port map( A => lpf_filter_inst_lpf_q_n1, Z
                           => lpf_filter_inst_lpf_q_n61);
   lpf_filter_inst_lpf_q_U45 : INVD1 port map( A => lpf_filter_inst_lpf_q_n2, Z
                           => lpf_filter_inst_lpf_q_n35);
   lpf_filter_inst_lpf_q_U44 : INVD1 port map( A => lpf_filter_inst_lpf_q_n2, Z
                           => lpf_filter_inst_lpf_q_n34);
   lpf_filter_inst_lpf_q_U43 : INVD1 port map( A => lpf_filter_inst_lpf_q_n2, Z
                           => lpf_filter_inst_lpf_q_n33);
   lpf_filter_inst_lpf_q_U42 : INVD1 port map( A => lpf_filter_inst_lpf_q_n2, Z
                           => lpf_filter_inst_lpf_q_n32);
   lpf_filter_inst_lpf_q_U41 : INVD1 port map( A => lpf_filter_inst_lpf_q_n2, Z
                           => lpf_filter_inst_lpf_q_n31);
   lpf_filter_inst_lpf_q_U40 : INVD1 port map( A => lpf_filter_inst_lpf_q_n2, Z
                           => lpf_filter_inst_lpf_q_n30);
   lpf_filter_inst_lpf_q_U39 : OAI21M20D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_12_port, 
                           A2 => lpf_filter_inst_lpf_q_n200, B => 
                           lpf_filter_inst_lpf_q_n199, Z => filter_out_q_0_port
                           );
   lpf_filter_inst_lpf_q_U38 : OAI21M20D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_13_port, 
                           A2 => lpf_filter_inst_lpf_q_n200, B => 
                           lpf_filter_inst_lpf_q_n199, Z => filter_out_q_1_port
                           );
   lpf_filter_inst_lpf_q_U37 : NAN4D1 port map( A1 => filter_out_q_4_port, A2 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_22_port, 
                           A3 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_21_port, 
                           A4 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_20_port, Z 
                           => lpf_filter_inst_lpf_q_n197);
   lpf_filter_inst_lpf_q_U36 : OAI21M20D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_15_port, 
                           A2 => lpf_filter_inst_lpf_q_n200, B => 
                           lpf_filter_inst_lpf_q_n199, Z => filter_out_q_3_port
                           );
   lpf_filter_inst_lpf_q_U35 : OAI21M20D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_14_port, 
                           A2 => lpf_filter_inst_lpf_q_n200, B => 
                           lpf_filter_inst_lpf_q_n199, Z => filter_out_q_2_port
                           );
   lpf_filter_inst_lpf_q_U34 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_sub_280_carry_18_port, Z => 
                           lpf_filter_inst_lpf_q_p141_1_19_port);
   lpf_filter_inst_lpf_q_U33 : NAN4D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_19_port, 
                           A2 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_18_port, 
                           A3 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_17_port, 
                           A4 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_16_port, Z 
                           => lpf_filter_inst_lpf_q_n198);
   lpf_filter_inst_lpf_q_U32 : INVD1 port map( A => lpf_filter_inst_lpf_q_n30, 
                           Z => lpf_filter_inst_lpf_q_n29);
   lpf_filter_inst_lpf_q_U31 : INVD1 port map( A => lpf_filter_inst_lpf_q_n30, 
                           Z => lpf_filter_inst_lpf_q_n4);
   lpf_filter_inst_lpf_q_U30 : INVD1 port map( A => lpf_filter_inst_lpf_q_n3, Z
                           => lpf_filter_inst_lpf_q_n5);
   lpf_filter_inst_lpf_q_U29 : INVD1 port map( A => lpf_filter_inst_lpf_q_n31, 
                           Z => lpf_filter_inst_lpf_q_n6);
   lpf_filter_inst_lpf_q_U28 : INVD1 port map( A => lpf_filter_inst_lpf_q_n35, 
                           Z => lpf_filter_inst_lpf_q_n7);
   lpf_filter_inst_lpf_q_U27 : INVD1 port map( A => lpf_filter_inst_lpf_q_n3, Z
                           => lpf_filter_inst_lpf_q_n8);
   lpf_filter_inst_lpf_q_U26 : INVD1 port map( A => lpf_filter_inst_lpf_q_n35, 
                           Z => lpf_filter_inst_lpf_q_n9);
   lpf_filter_inst_lpf_q_U25 : INVD1 port map( A => lpf_filter_inst_lpf_q_n35, 
                           Z => lpf_filter_inst_lpf_q_n10);
   lpf_filter_inst_lpf_q_U24 : INVD1 port map( A => lpf_filter_inst_lpf_q_n35, 
                           Z => lpf_filter_inst_lpf_q_n11);
   lpf_filter_inst_lpf_q_U23 : INVD1 port map( A => lpf_filter_inst_lpf_q_n34, 
                           Z => lpf_filter_inst_lpf_q_n12);
   lpf_filter_inst_lpf_q_U22 : INVD1 port map( A => lpf_filter_inst_lpf_q_n33, 
                           Z => lpf_filter_inst_lpf_q_n13);
   lpf_filter_inst_lpf_q_U21 : INVD1 port map( A => lpf_filter_inst_lpf_q_n32, 
                           Z => lpf_filter_inst_lpf_q_n14);
   lpf_filter_inst_lpf_q_U20 : INVD1 port map( A => lpf_filter_inst_lpf_q_n34, 
                           Z => lpf_filter_inst_lpf_q_n15);
   lpf_filter_inst_lpf_q_U15 : INVD1 port map( A => lpf_filter_inst_lpf_q_n34, 
                           Z => lpf_filter_inst_lpf_q_n16);
   lpf_filter_inst_lpf_q_U14 : INVD1 port map( A => lpf_filter_inst_lpf_q_n34, 
                           Z => lpf_filter_inst_lpf_q_n17);
   lpf_filter_inst_lpf_q_U13 : INVD1 port map( A => lpf_filter_inst_lpf_q_n33, 
                           Z => lpf_filter_inst_lpf_q_n18);
   lpf_filter_inst_lpf_q_U12 : INVD1 port map( A => lpf_filter_inst_lpf_q_n33, 
                           Z => lpf_filter_inst_lpf_q_n19);
   lpf_filter_inst_lpf_q_U11 : INVD1 port map( A => lpf_filter_inst_lpf_q_n33, 
                           Z => lpf_filter_inst_lpf_q_n20);
   lpf_filter_inst_lpf_q_U10 : INVD1 port map( A => lpf_filter_inst_lpf_q_n32, 
                           Z => lpf_filter_inst_lpf_q_n21);
   lpf_filter_inst_lpf_q_U9 : INVD1 port map( A => lpf_filter_inst_lpf_q_n32, Z
                           => lpf_filter_inst_lpf_q_n22);
   lpf_filter_inst_lpf_q_U8 : INVD1 port map( A => lpf_filter_inst_lpf_q_n32, Z
                           => lpf_filter_inst_lpf_q_n23);
   lpf_filter_inst_lpf_q_U7 : INVD1 port map( A => lpf_filter_inst_lpf_q_n31, Z
                           => lpf_filter_inst_lpf_q_n24);
   lpf_filter_inst_lpf_q_U6 : INVD1 port map( A => lpf_filter_inst_lpf_q_n31, Z
                           => lpf_filter_inst_lpf_q_n25);
   lpf_filter_inst_lpf_q_U5 : INVD1 port map( A => lpf_filter_inst_lpf_q_n31, Z
                           => lpf_filter_inst_lpf_q_n26);
   lpf_filter_inst_lpf_q_U4 : INVD1 port map( A => lpf_filter_inst_lpf_q_n30, Z
                           => lpf_filter_inst_lpf_q_n27);
   lpf_filter_inst_lpf_q_U3 : INVD1 port map( A => lpf_filter_inst_lpf_q_n30, Z
                           => lpf_filter_inst_lpf_q_n28);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_36_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_24_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_37_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_25_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_38_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_26_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_39_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_27_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_40_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_28_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_41_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_29_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_42_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_30_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_43_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_31_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_44_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_32_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_45_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_33_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_46_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_34_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_25_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_47_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_35_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_84_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_72_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_85_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_73_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_86_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_74_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_87_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_75_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_88_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_76_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_89_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_77_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_90_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_78_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_91_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_79_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_92_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_80_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_93_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_81_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_94_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_82_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_21_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_95_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_83_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_132_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_120_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_133_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_121_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_134_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_122_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_135_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_123_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_136_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_124_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_137_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_125_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_138_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_126_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_139_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_127_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_140_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_128_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_141_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_129_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_142_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_130_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_17_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_143_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_131_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_227_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_215_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_228_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_216_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_229_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_217_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_230_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_218_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_231_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_219_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_232_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_220_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_233_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_221_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_234_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_222_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_235_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_223_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_236_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_224_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_237_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_225_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_9_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_238_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_226_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_275_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_263_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_276_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_264_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_277_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_265_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_278_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_266_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_279_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_267_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_280_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_268_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_281_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_269_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_282_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_270_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_283_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_271_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_284_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_272_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_285_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_273_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_5_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_286_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_274_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_323_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_311_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_324_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_312_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_325_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_313_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_326_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_314_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_327_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_315_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_328_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_316_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_329_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_317_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_330_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_318_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_331_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_319_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_332_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_320_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_333_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_321_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_1_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_334_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_322_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_190_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_178_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_179_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_t11_14_0_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_181_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_169_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_182_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_170_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_183_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_171_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_184_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_172_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_185_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_173_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_186_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_174_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_187_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_175_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_188_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_176_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_189_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_177_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_13_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_180_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_168_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_202_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_190_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_214_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_202_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_226_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_214_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_250_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_238_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_262_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_250_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_274_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_262_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_298_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_286_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_310_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_298_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_322_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_310_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_11 : DFFRPQ1 port map( D => 
                           mixer_out_q_11_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_334_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_35_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_23_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_59_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_47_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_71_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_59_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_83_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_71_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_107_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_95_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_119_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_107_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_131_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_119_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_155_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_143_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_167_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_155_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_p232_2_17, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n16, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_167_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_24_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_12_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_48_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n27, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_36_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_60_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_48_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_72_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_60_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_96_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_84_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_108_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_96_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_120_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_108_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_144_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_132_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_156_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_144_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_t11_14_0_port, CK => clk, RB 
                           => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_156_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_192_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_180_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_193_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_181_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_194_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_182_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_195_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_183_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_196_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_184_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_197_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_185_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_198_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_186_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_199_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_187_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_200_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_188_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_201_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_189_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_204_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_192_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_205_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_193_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_206_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_194_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_207_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_195_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_208_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_196_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_209_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_197_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_210_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_198_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_211_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_199_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_212_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_200_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_213_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_201_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_216_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_204_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_217_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_205_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_218_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_206_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_219_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_207_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_220_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_208_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_221_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_209_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_222_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_210_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_223_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_211_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_224_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_212_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_225_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n13, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_213_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_240_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_228_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_241_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_229_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_242_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_230_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_243_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_231_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_244_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_232_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_245_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_233_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_246_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_234_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_247_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_235_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_248_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_236_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_249_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_237_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_252_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_240_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_253_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_241_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_254_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_242_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_255_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_243_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_256_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_244_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_257_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_245_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_258_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_246_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_259_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_247_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_260_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_248_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_261_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_249_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_264_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_252_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_265_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_253_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_266_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_254_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_267_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_255_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_268_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_256_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_269_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_257_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_270_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_258_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_271_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_259_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_272_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_260_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_273_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n9, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_261_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_288_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_276_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_289_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_277_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_290_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_278_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_291_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_279_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_292_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_280_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_293_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_281_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_294_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_282_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_295_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_283_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_296_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_284_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_297_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_285_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_300_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_288_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_301_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_289_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_302_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_290_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_303_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_291_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_304_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_292_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_305_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_293_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_306_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_294_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_307_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_295_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_308_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_296_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_309_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_297_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_312_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_300_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_313_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_301_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_314_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_302_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_315_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_303_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_316_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_304_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_317_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_305_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_318_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_306_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_319_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_307_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_320_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_308_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_321_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n5, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_309_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_1 : DFFRPQ1 port map( D => 
                           mixer_out_q_1_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_324_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_2 : DFFRPQ1 port map( D => 
                           mixer_out_q_2_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_325_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_3 : DFFRPQ1 port map( D => 
                           mixer_out_q_3_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_326_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_4 : DFFRPQ1 port map( D => 
                           mixer_out_q_4_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_327_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_5 : DFFRPQ1 port map( D => 
                           mixer_out_q_5_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_328_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_6 : DFFRPQ1 port map( D => 
                           mixer_out_q_6_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_329_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_7 : DFFRPQ1 port map( D => 
                           mixer_out_q_7_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_330_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_8 : DFFRPQ1 port map( D => 
                           mixer_out_q_8_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_331_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_9 : DFFRPQ1 port map( D => 
                           mixer_out_q_9_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_332_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_10 : DFFRPQ1 port map( D => 
                           mixer_out_q_10_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_333_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_25_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_13_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_26_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_14_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_27_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_15_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_28_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_16_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_29_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_17_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_30_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_18_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_31_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_19_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_32_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_20_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_33_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_21_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_26_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_34_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_22_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_49_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_37_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_50_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_38_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_51_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_39_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_52_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_40_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_53_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_41_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_54_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_42_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_55_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_43_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_56_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_44_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_57_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_45_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_24_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_58_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_46_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_61_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n26, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_49_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_62_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_50_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_63_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_51_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_64_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_52_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_65_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_53_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_66_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_54_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_67_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_55_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_68_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_56_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_69_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_57_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_23_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_70_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_58_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_73_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_61_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_74_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n25, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_62_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_75_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_63_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_76_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_64_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_77_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_65_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_78_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_66_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_79_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_67_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_80_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_68_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_81_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_69_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_22_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_82_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n24, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_70_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_97_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_85_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_98_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_86_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_99_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_87_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_100_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n23, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_88_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_101_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_89_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_102_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_90_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_103_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_91_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_104_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_92_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_105_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_93_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_20_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_106_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_94_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_109_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_97_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_110_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_98_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_111_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_99_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_112_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_100_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_113_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n22, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_101_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_114_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_102_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_115_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_103_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_116_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_104_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_117_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_105_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_19_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_118_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_106_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_121_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_109_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_122_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_110_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_123_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_111_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_124_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_112_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_125_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_113_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_126_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n21, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_114_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_127_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_115_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_128_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_116_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_129_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_117_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_18_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_130_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n20, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_118_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_145_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_133_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_146_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_134_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_147_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_135_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_148_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_136_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_149_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_137_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_150_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_138_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_151_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_139_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_152_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n19, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_140_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_153_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_141_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_16_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_154_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_142_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_157_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_145_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_158_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_146_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_159_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_147_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_160_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_148_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_161_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_149_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_162_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_150_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_163_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_151_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_164_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_152_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_165_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n18, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_153_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_15_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_166_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_154_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_168_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_157_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_169_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_158_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_170_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_159_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_171_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_160_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_172_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_161_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_173_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_162_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_174_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_163_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_175_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_164_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_176_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_165_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_14_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_177_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n17, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_166_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_12_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_191_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_179_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_11_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_203_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n15, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_191_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_10_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_215_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n14, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_203_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_8_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_239_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n12, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_227_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_7_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_251_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n11, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_239_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_6_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_263_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n10, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_251_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_4_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_287_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n8, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_275_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_3_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_299_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n7, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_287_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_2_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_311_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n6, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_299_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_0_0 : DFFRPQ1 port map( D => 
                           mixer_out_q_0_port, CK => clk, RB => 
                           lpf_filter_inst_lpf_q_n4, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_323_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_11 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_23_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n28, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_11_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_0 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_12_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_0_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_1 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_13_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_1_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_2 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_14_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_2_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_3 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_15_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_3_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_4 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_16_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_4_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_5 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_17_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_5_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_6 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_18_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_6_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_7 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_19_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_7_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_8 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_20_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_8_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_9 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_21_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_9_port);
   lpf_filter_inst_lpf_q_arx_input_reg_reg_27_10 : DFFRPQ1 port map( D => 
                           lpf_filter_inst_lpf_q_arx_input_reg_22_port, CK => 
                           clk, RB => lpf_filter_inst_lpf_q_n29, Q => 
                           lpf_filter_inst_lpf_q_arx_input_reg_10_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_20 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_19, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_20_port, 
                           CO => lpf_filter_inst_lpf_q_n_1371, S => 
                           lpf_filter_inst_lpf_q_p206_3_20_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_19, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_20_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_19_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_18, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_19_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_18_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_17, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_17_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_16, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_16_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_15, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_15_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_14, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_14_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_13, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_13_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_12, B => 
                           lpf_filter_inst_lpf_q_n48, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_12_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_11, B => 
                           lpf_filter_inst_lpf_q_n47, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_11_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_10, B => 
                           lpf_filter_inst_lpf_q_n46, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_10_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_9, B => 
                           lpf_filter_inst_lpf_q_n45, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_9_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_8, B => 
                           lpf_filter_inst_lpf_q_n44, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_8_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_7, B => 
                           lpf_filter_inst_lpf_q_n43, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_7_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_6, B => 
                           lpf_filter_inst_lpf_q_n42, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_6_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_5, B => 
                           lpf_filter_inst_lpf_q_n41, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_5_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_4, B => 
                           lpf_filter_inst_lpf_q_n40, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_4_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_285_U2_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_3, B => 
                           lpf_filter_inst_lpf_q_n39, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_285_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_p206_3_3_port);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_17, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_177_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_11, 
                           CO => lpf_filter_inst_lpf_q_p232_2_12, S => 
                           lpf_filter_inst_lpf_q_p232_2_11);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_177_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_176_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_10, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_11, S
                           => lpf_filter_inst_lpf_q_p232_2_10);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_176_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_175_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_9, CO
                           => lpf_filter_inst_lpf_q_add_1_root_add_286_carry_10
                           , S => lpf_filter_inst_lpf_q_p232_2_9);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_175_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_174_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_8, CO
                           => lpf_filter_inst_lpf_q_add_1_root_add_286_carry_9,
                           S => lpf_filter_inst_lpf_q_p232_2_8);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_174_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_173_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_7, CO
                           => lpf_filter_inst_lpf_q_add_1_root_add_286_carry_8,
                           S => lpf_filter_inst_lpf_q_p232_2_7);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_173_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_172_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_6, CO
                           => lpf_filter_inst_lpf_q_add_1_root_add_286_carry_7,
                           S => lpf_filter_inst_lpf_q_p232_2_6);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_172_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_171_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_5, CO
                           => lpf_filter_inst_lpf_q_add_1_root_add_286_carry_6,
                           S => lpf_filter_inst_lpf_q_p232_2_5);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_171_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_170_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_4, CO
                           => lpf_filter_inst_lpf_q_add_1_root_add_286_carry_5,
                           S => lpf_filter_inst_lpf_q_p232_2_4);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_170_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_169_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_3, CO
                           => lpf_filter_inst_lpf_q_add_1_root_add_286_carry_4,
                           S => lpf_filter_inst_lpf_q_p232_2_3);
   lpf_filter_inst_lpf_q_add_1_root_add_286_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_169_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_168_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_286_carry_2, CO
                           => lpf_filter_inst_lpf_q_add_1_root_add_286_carry_3,
                           S => lpf_filter_inst_lpf_q_p232_2_2);
   lpf_filter_inst_lpf_q_sub_280_U2_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_11_port, B => 
                           lpf_filter_inst_lpf_q_n61, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_17_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_18_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_17_port);
   lpf_filter_inst_lpf_q_sub_280_U2_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_10_port, B => 
                           lpf_filter_inst_lpf_q_n61, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_16_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_17_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_16_port);
   lpf_filter_inst_lpf_q_sub_280_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_9_port, B => 
                           lpf_filter_inst_lpf_q_n61, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_15_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_16_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_15_port);
   lpf_filter_inst_lpf_q_sub_280_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_8_port, B => 
                           lpf_filter_inst_lpf_q_n61, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_14_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_15_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_14_port);
   lpf_filter_inst_lpf_q_sub_280_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_7_port, B => 
                           lpf_filter_inst_lpf_q_n61, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_13_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_14_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_13_port);
   lpf_filter_inst_lpf_q_sub_280_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_6_port, B => 
                           lpf_filter_inst_lpf_q_n61, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_12_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_13_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_12_port);
   lpf_filter_inst_lpf_q_sub_280_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_5_port, B => 
                           lpf_filter_inst_lpf_q_n60, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_11_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_12_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_11_port);
   lpf_filter_inst_lpf_q_sub_280_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_4_port, B => 
                           lpf_filter_inst_lpf_q_n59, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_10_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_11_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_10_port);
   lpf_filter_inst_lpf_q_sub_280_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_3_port, B => 
                           lpf_filter_inst_lpf_q_n58, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_9_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_10_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_9_port);
   lpf_filter_inst_lpf_q_sub_280_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_2_port, B => 
                           lpf_filter_inst_lpf_q_n57, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_8_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_9_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_8_port);
   lpf_filter_inst_lpf_q_sub_280_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_1_port, B => 
                           lpf_filter_inst_lpf_q_n56, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_7_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_8_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_7_port);
   lpf_filter_inst_lpf_q_sub_280_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n117, B => 
                           lpf_filter_inst_lpf_q_n55, CI => 
                           lpf_filter_inst_lpf_q_sub_280_carry_6_port, CO => 
                           lpf_filter_inst_lpf_q_sub_280_carry_7_port, S => 
                           lpf_filter_inst_lpf_q_p141_1_6_port);
   lpf_filter_inst_lpf_q_add_284_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_11_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_15_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_13, CO => 
                           lpf_filter_inst_lpf_q_p206_2_14_port, S => 
                           lpf_filter_inst_lpf_q_p206_2_13_port);
   lpf_filter_inst_lpf_q_add_284_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_10_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_15_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_12, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_13, S => 
                           lpf_filter_inst_lpf_q_p206_2_12_port);
   lpf_filter_inst_lpf_q_add_284_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_9_port, B => 
                           lpf_filter_inst_lpf_q_pair13_15_11_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_11, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_12, S => 
                           lpf_filter_inst_lpf_q_p206_2_11_port);
   lpf_filter_inst_lpf_q_add_284_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_8_port, B => 
                           lpf_filter_inst_lpf_q_pair13_15_10_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_10, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_11, S => 
                           lpf_filter_inst_lpf_q_p206_2_10_port);
   lpf_filter_inst_lpf_q_add_284_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_7_port, B => 
                           lpf_filter_inst_lpf_q_pair13_15_9_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_9, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_10, S => 
                           lpf_filter_inst_lpf_q_p206_2_9_port);
   lpf_filter_inst_lpf_q_add_284_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_6_port, B => 
                           lpf_filter_inst_lpf_q_pair13_15_8_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_8, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_9, S => 
                           lpf_filter_inst_lpf_q_p206_2_8_port);
   lpf_filter_inst_lpf_q_add_284_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_5_port, B => 
                           lpf_filter_inst_lpf_q_pair13_15_7_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_7, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_8, S => 
                           lpf_filter_inst_lpf_q_p206_2_7_port);
   lpf_filter_inst_lpf_q_add_284_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_4_port, B => 
                           lpf_filter_inst_lpf_q_pair13_15_6_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_6, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_7, S => 
                           lpf_filter_inst_lpf_q_p206_2_6_port);
   lpf_filter_inst_lpf_q_add_284_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_3_port, B => 
                           lpf_filter_inst_lpf_q_pair13_15_5_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_5, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_6, S => 
                           lpf_filter_inst_lpf_q_p206_2_5_port);
   lpf_filter_inst_lpf_q_add_284_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_2_port, B => 
                           lpf_filter_inst_lpf_q_pair13_15_4_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_4, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_5, S => 
                           lpf_filter_inst_lpf_q_p206_2_4_port);
   lpf_filter_inst_lpf_q_add_284_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_4, B => 
                           lpf_filter_inst_lpf_q_pair13_15_3_port, CI => 
                           lpf_filter_inst_lpf_q_add_284_carry_3, CO => 
                           lpf_filter_inst_lpf_q_add_284_carry_4, S => 
                           lpf_filter_inst_lpf_q_p206_2_3_port);
   lpf_filter_inst_lpf_q_U19 : OR4D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_20_port, 
                           A2 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_21_port, 
                           A3 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_22_port, 
                           A4 => filter_out_q_4_port, Z => 
                           lpf_filter_inst_lpf_q_n196);
   lpf_filter_inst_lpf_q_U18 : OR4D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_16_port, 
                           A2 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_17_port, 
                           A3 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_18_port, 
                           A4 => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_19_port, Z 
                           => lpf_filter_inst_lpf_q_n195);
   lpf_filter_inst_lpf_q_U17 : OAI22D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_n198, A2 => 
                           lpf_filter_inst_lpf_q_n197, B1 => 
                           lpf_filter_inst_lpf_q_n196, B2 => 
                           lpf_filter_inst_lpf_q_n195, Z => 
                           lpf_filter_inst_lpf_q_n200);
   lpf_filter_inst_lpf_q_U16 : OR2D1 port map( A1 => lpf_filter_inst_lpf_q_n200
                           , A2 => filter_out_q_4_port, Z => 
                           lpf_filter_inst_lpf_q_n199);
   lpf_filter_inst_lpf_q_add_273_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_156_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_179_port, Z => 
                           lpf_filter_inst_lpf_q_p206_1_3);
   lpf_filter_inst_lpf_q_add_273_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_156_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_179_port, Z => 
                           lpf_filter_inst_lpf_q_add_273_n1);
   lpf_filter_inst_lpf_q_add_273_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_180_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_157_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_n1, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_2_port, S => 
                           lpf_filter_inst_lpf_q_p206_1_4);
   lpf_filter_inst_lpf_q_add_273_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_181_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_158_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_2_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_3_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_2_port);
   lpf_filter_inst_lpf_q_add_273_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_182_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_159_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_3_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_4_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_3_port);
   lpf_filter_inst_lpf_q_add_273_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_183_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_160_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_4_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_5_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_4_port);
   lpf_filter_inst_lpf_q_add_273_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_184_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_161_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_5_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_6_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_5_port);
   lpf_filter_inst_lpf_q_add_273_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_185_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_162_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_6_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_7_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_6_port);
   lpf_filter_inst_lpf_q_add_273_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_186_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_163_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_7_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_8_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_7_port);
   lpf_filter_inst_lpf_q_add_273_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_187_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_164_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_8_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_9_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_8_port);
   lpf_filter_inst_lpf_q_add_273_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_188_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_165_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_9_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_10_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_9_port);
   lpf_filter_inst_lpf_q_add_273_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_189_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_166_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_10_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_11_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_10_port);
   lpf_filter_inst_lpf_q_add_273_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_190_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_167_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_11_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_carry_12_port, S => 
                           lpf_filter_inst_lpf_q_pair13_15_11_port);
   lpf_filter_inst_lpf_q_add_273_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_190_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_167_port, CI => 
                           lpf_filter_inst_lpf_q_add_273_carry_12_port, CO => 
                           lpf_filter_inst_lpf_q_add_273_n_1321, S => 
                           lpf_filter_inst_lpf_q_p206_2_15_port);
   lpf_filter_inst_lpf_q_add_272_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_144_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_191_port, Z => 
                           lpf_filter_inst_lpf_q_n117);
   lpf_filter_inst_lpf_q_add_272_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_144_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_191_port, Z => 
                           lpf_filter_inst_lpf_q_add_272_n1);
   lpf_filter_inst_lpf_q_add_272_U1_12 : EXOR3D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_202_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_155_port, A3 => 
                           lpf_filter_inst_lpf_q_add_272_carry_12_port, Z => 
                           lpf_filter_inst_lpf_q_pair12_16_12_port);
   lpf_filter_inst_lpf_q_add_272_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_192_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_145_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_n1, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_2_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_1_port);
   lpf_filter_inst_lpf_q_add_272_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_193_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_146_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_2_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_3_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_2_port);
   lpf_filter_inst_lpf_q_add_272_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_194_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_147_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_3_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_4_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_3_port);
   lpf_filter_inst_lpf_q_add_272_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_195_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_148_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_4_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_5_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_4_port);
   lpf_filter_inst_lpf_q_add_272_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_196_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_149_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_5_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_6_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_5_port);
   lpf_filter_inst_lpf_q_add_272_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_197_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_150_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_6_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_7_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_6_port);
   lpf_filter_inst_lpf_q_add_272_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_198_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_151_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_7_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_8_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_7_port);
   lpf_filter_inst_lpf_q_add_272_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_199_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_152_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_8_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_9_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_8_port);
   lpf_filter_inst_lpf_q_add_272_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_200_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_153_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_9_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_10_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_9_port);
   lpf_filter_inst_lpf_q_add_272_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_201_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_154_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_10_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_11_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_10_port);
   lpf_filter_inst_lpf_q_add_272_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_202_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_155_port, CI => 
                           lpf_filter_inst_lpf_q_add_272_carry_11_port, CO => 
                           lpf_filter_inst_lpf_q_add_272_carry_12_port, S => 
                           lpf_filter_inst_lpf_q_pair12_16_11_port);
   lpf_filter_inst_lpf_q_add_271_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_132_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_203_port, Z => 
                           lpf_filter_inst_lpf_q_n74);
   lpf_filter_inst_lpf_q_add_271_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_132_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_203_port, Z => 
                           lpf_filter_inst_lpf_q_add_271_n1);
   lpf_filter_inst_lpf_q_add_271_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_204_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_133_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_n1, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_2_port, S => 
                           lpf_filter_inst_lpf_q_n67);
   lpf_filter_inst_lpf_q_add_271_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_205_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_134_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_2_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_3_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_2_port);
   lpf_filter_inst_lpf_q_add_271_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_206_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_135_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_3_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_4_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_3_port);
   lpf_filter_inst_lpf_q_add_271_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_207_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_136_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_4_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_5_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_4_port);
   lpf_filter_inst_lpf_q_add_271_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_208_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_137_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_5_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_6_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_5_port);
   lpf_filter_inst_lpf_q_add_271_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_209_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_138_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_6_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_7_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_6_port);
   lpf_filter_inst_lpf_q_add_271_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_210_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_139_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_7_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_8_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_7_port);
   lpf_filter_inst_lpf_q_add_271_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_211_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_140_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_8_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_9_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_8_port);
   lpf_filter_inst_lpf_q_add_271_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_212_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_141_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_9_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_10_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_9_port);
   lpf_filter_inst_lpf_q_add_271_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_213_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_142_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_10_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_11_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_10_port);
   lpf_filter_inst_lpf_q_add_271_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_214_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_143_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_11_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_carry_12_port, S => 
                           lpf_filter_inst_lpf_q_pair11_17_11_port);
   lpf_filter_inst_lpf_q_add_271_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_214_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_143_port, CI => 
                           lpf_filter_inst_lpf_q_add_271_carry_12_port, CO => 
                           lpf_filter_inst_lpf_q_add_271_n_1316, S => 
                           lpf_filter_inst_lpf_q_pair11_17_12_port);
   lpf_filter_inst_lpf_q_add_268_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_84_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_251_port, Z => 
                           lpf_filter_inst_lpf_q_pair7_21_0_port);
   lpf_filter_inst_lpf_q_add_268_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_84_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_251_port, Z => 
                           lpf_filter_inst_lpf_q_add_268_n1);
   lpf_filter_inst_lpf_q_add_268_U1_12 : EXOR3D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_262_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_95_port, A3 => 
                           lpf_filter_inst_lpf_q_add_268_carry_12_port, Z => 
                           lpf_filter_inst_lpf_q_pair7_21_12_port);
   lpf_filter_inst_lpf_q_add_268_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_252_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_85_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_n1, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_2_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_1_port);
   lpf_filter_inst_lpf_q_add_268_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_253_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_86_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_2_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_3_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_2_port);
   lpf_filter_inst_lpf_q_add_268_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_254_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_87_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_3_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_4_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_3_port);
   lpf_filter_inst_lpf_q_add_268_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_255_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_88_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_4_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_5_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_4_port);
   lpf_filter_inst_lpf_q_add_268_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_256_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_89_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_5_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_6_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_5_port);
   lpf_filter_inst_lpf_q_add_268_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_257_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_90_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_6_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_7_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_6_port);
   lpf_filter_inst_lpf_q_add_268_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_258_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_91_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_7_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_8_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_7_port);
   lpf_filter_inst_lpf_q_add_268_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_259_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_92_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_8_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_9_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_8_port);
   lpf_filter_inst_lpf_q_add_268_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_260_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_93_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_9_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_10_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_9_port);
   lpf_filter_inst_lpf_q_add_268_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_261_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_94_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_10_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_11_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_10_port);
   lpf_filter_inst_lpf_q_add_268_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_262_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_95_port, CI => 
                           lpf_filter_inst_lpf_q_add_268_carry_11_port, CO => 
                           lpf_filter_inst_lpf_q_add_268_carry_12_port, S => 
                           lpf_filter_inst_lpf_q_pair7_21_11_port);
   lpf_filter_inst_lpf_q_add_264_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_12_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_323_port, Z => 
                           lpf_filter_inst_lpf_q_pair1_27_0_port);
   lpf_filter_inst_lpf_q_add_264_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_12_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_323_port, Z => 
                           lpf_filter_inst_lpf_q_add_264_n1);
   lpf_filter_inst_lpf_q_add_264_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_324_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_13_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_n1, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_2_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_1_port);
   lpf_filter_inst_lpf_q_add_264_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_325_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_14_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_2_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_3_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_2_port);
   lpf_filter_inst_lpf_q_add_264_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_326_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_15_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_3_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_4_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_3_port);
   lpf_filter_inst_lpf_q_add_264_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_327_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_16_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_4_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_5_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_4_port);
   lpf_filter_inst_lpf_q_add_264_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_328_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_17_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_5_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_6_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_5_port);
   lpf_filter_inst_lpf_q_add_264_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_329_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_18_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_6_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_7_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_6_port);
   lpf_filter_inst_lpf_q_add_264_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_330_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_19_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_7_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_8_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_7_port);
   lpf_filter_inst_lpf_q_add_264_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_331_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_20_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_8_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_9_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_8_port);
   lpf_filter_inst_lpf_q_add_264_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_332_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_21_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_9_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_10_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_9_port);
   lpf_filter_inst_lpf_q_add_264_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_333_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_22_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_10_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_11_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_10_port);
   lpf_filter_inst_lpf_q_add_264_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_334_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_23_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_11_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_carry_12_port, S => 
                           lpf_filter_inst_lpf_q_pair1_27_11_port);
   lpf_filter_inst_lpf_q_add_264_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_334_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_23_port, CI => 
                           lpf_filter_inst_lpf_q_add_264_carry_12_port, CO => 
                           lpf_filter_inst_lpf_q_add_264_n_1311, S => 
                           lpf_filter_inst_lpf_q_pair1_27_12_port);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_0_port, A2 => 
                           mixer_out_q_0_port, Z => 
                           lpf_filter_inst_lpf_q_pair0_28_0);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_0_port, A2 => 
                           mixer_out_q_0_port, Z => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_n1);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_12 : EXOR3D1 port map( A1 => 
                           mixer_out_q_11_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_11_port, A3 => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_12_port, Z 
                           => lpf_filter_inst_lpf_q_pair0_28_12);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_1 : ADFULD1 port map( A => 
                           mixer_out_q_1_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_1_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_2_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_1);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_2 : ADFULD1 port map( A => 
                           mixer_out_q_2_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_2_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_2);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_3 : ADFULD1 port map( A => 
                           mixer_out_q_3_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_3_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_3);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_4 : ADFULD1 port map( A => 
                           mixer_out_q_4_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_4_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_4);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_5 : ADFULD1 port map( A => 
                           mixer_out_q_5_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_5_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_5);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_6 : ADFULD1 port map( A => 
                           mixer_out_q_6_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_6_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_6);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_7 : ADFULD1 port map( A => 
                           mixer_out_q_7_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_7_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_7);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_8 : ADFULD1 port map( A => 
                           mixer_out_q_8_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_8_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_8);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_9 : ADFULD1 port map( A => 
                           mixer_out_q_9_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_9_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_9);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_10 : ADFULD1 port map( A => 
                           mixer_out_q_10_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_10_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_10);
   lpf_filter_inst_lpf_q_add_5_root_add_292_U1_11 : ADFULD1 port map( A => 
                           mixer_out_q_11_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_11_port, CI => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_5_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_pair0_28_11);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair12_16_1_port, A2 => 
                           lpf_filter_inst_lpf_q_pair1_27_0_port, Z => 
                           lpf_filter_inst_lpf_q_t0_1_1);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair12_16_1_port, A2 => 
                           lpf_filter_inst_lpf_q_pair1_27_0_port, Z => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_n1);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_14 : EXOR3D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair1_27_12_port, A2 => 
                           lpf_filter_inst_lpf_q_n1, A3 => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_14_port, Z 
                           => lpf_filter_inst_lpf_q_t0_1_14);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_1_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_2_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_2);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_2_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_3_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_3);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_3_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_4_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_4);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_4_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_5_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_5);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_5_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_6_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_6);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_6_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_7_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_7);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_7_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_8_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_8);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_8_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_9_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_9);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_9_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_10_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_10);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_10_port, B => 
                           lpf_filter_inst_lpf_q_pair12_16_11_port, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_11);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_11_port, B => 
                           lpf_filter_inst_lpf_q_n1, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_12);
   lpf_filter_inst_lpf_q_add_4_root_add_292_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair1_27_12_port, B => 
                           lpf_filter_inst_lpf_q_n1, CI => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_4_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_t0_1_13);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_p141_1_2_port, A2 => 
                           lpf_filter_inst_lpf_q_t11_14_0_port, Z => 
                           lpf_filter_inst_lpf_q_n156);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_p141_1_2_port, A2 => 
                           lpf_filter_inst_lpf_q_t11_14_0_port, Z => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_n1);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_1_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_3_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_n155);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_2_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_4_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_n154);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_3_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_5_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_n153);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_4_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_6_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_n152);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_5_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_7_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_n151);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_6_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_8_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_n150);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_7_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_9_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_n149);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_8_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_10_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_n148);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_9_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_11_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_n147);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_10_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_12_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_n146);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_11_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_13_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_n145);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_12_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_14_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_n144);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_13_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_15_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_n143);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_14_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_16_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_n142);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_15_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_17_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_q_n141);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_16_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_19_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_q_n140);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_20 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_17_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_19_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_q_n139);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_21 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_18_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_19_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_q_n138);
   lpf_filter_inst_lpf_q_add_7_root_add_292_U1_22 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_18_port, B => 
                           lpf_filter_inst_lpf_q_p141_1_19_port, CI => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_7_root_add_292_n_1079, S 
                           => lpf_filter_inst_lpf_q_n137);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_3_port, A2 => 
                           lpf_filter_inst_lpf_q_t3_7_1_port, Z => 
                           lpf_filter_inst_lpf_q_n135);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_3_port, A2 => 
                           lpf_filter_inst_lpf_q_t3_7_1_port, Z => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_n1);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_2_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_4_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_n134);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_3_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_5_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_n133);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_4_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_6_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_n132);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_5_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_7_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_n131);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_6_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_8_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_n130);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_7_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_9_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_n129);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_8_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_10_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_n128);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_9_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_11_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_n127);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_10_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_12_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_n126);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_11_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_13_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_n125);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_12_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_14_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_n124);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_13_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_15_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_n123);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_14_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_16_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_n122);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_15_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_17_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_n121);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_15_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_18_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_q_n120);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_15_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_19_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_q_n119);
   lpf_filter_inst_lpf_q_add_8_root_add_292_U1_20 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t3_7_15_port, B => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_19_port, CI => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_8_root_add_292_n_1089, S 
                           => lpf_filter_inst_lpf_q_n118);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_p206_3_3_port, A2 => 
                           lpf_filter_inst_lpf_q_n117, Z => 
                           lpf_filter_inst_lpf_q_t12_13_4);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_p206_3_3_port, A2 => 
                           lpf_filter_inst_lpf_q_n117, Z => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_n1);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_1_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_4_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_n1, CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_5);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_2_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_5_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_6);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_3_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_6_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_7);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_4_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_7_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_8);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_5_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_8_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_9);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_6_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_9_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_10);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_7_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_10_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_11);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_8_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_11_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_12);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_9_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_12_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_13);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_10_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_13_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_14);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair12_16_11_port, B => 
                           lpf_filter_inst_lpf_q_p206_3_14_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_15);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n1, B => 
                           lpf_filter_inst_lpf_q_p206_3_15_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_16);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n1, B => 
                           lpf_filter_inst_lpf_q_p206_3_16_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_17);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n1, B => 
                           lpf_filter_inst_lpf_q_p206_3_17_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_18);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n1, B => 
                           lpf_filter_inst_lpf_q_p206_3_18_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_19);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_20 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n1, B => 
                           lpf_filter_inst_lpf_q_p206_3_19_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_20);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_21 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n1, B => 
                           lpf_filter_inst_lpf_q_p206_3_20_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_q_t12_13_21);
   lpf_filter_inst_lpf_q_add_6_root_add_292_U1_22 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n1, B => 
                           lpf_filter_inst_lpf_q_p206_3_20_port, CI => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_6_root_add_292_n_1098, S 
                           => lpf_filter_inst_lpf_q_t12_13_22);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U2 : EXOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_q_n117, A2 => 
                           lpf_filter_inst_lpf_q_p206_1_3, Z => 
                           lpf_filter_inst_lpf_q_n181);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1 : AND2D1 port map( A1
                           => lpf_filter_inst_lpf_q_n117, A2 => 
                           lpf_filter_inst_lpf_q_p206_1_3, Z => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_n1);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_2 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_t12_13_2, B => 
                           lpf_filter_inst_lpf_q_n157, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_n1, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_n180);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_3 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_t12_13_3, B => 
                           lpf_filter_inst_lpf_q_n156, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_n179);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_4 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_t12_13_4, B => 
                           lpf_filter_inst_lpf_q_n155, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_n178);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_5 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_t12_13_5, B => 
                           lpf_filter_inst_lpf_q_n154, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_n177);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_6 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_t12_13_6, B => 
                           lpf_filter_inst_lpf_q_n153, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_n176);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_7 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_t12_13_7, B => 
                           lpf_filter_inst_lpf_q_n152, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_n175);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_8 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_t12_13_8, B => 
                           lpf_filter_inst_lpf_q_n151, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_n174);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_9 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_t12_13_9, B => 
                           lpf_filter_inst_lpf_q_n150, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_n173);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_10 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_10, B => 
                           lpf_filter_inst_lpf_q_n149, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_n172);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_11 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_11, B => 
                           lpf_filter_inst_lpf_q_n148, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_n171);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_12 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_12, B => 
                           lpf_filter_inst_lpf_q_n147, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_n170);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_13 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_13, B => 
                           lpf_filter_inst_lpf_q_n146, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_n169);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_14 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_14, B => 
                           lpf_filter_inst_lpf_q_n145, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_n168);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_15 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_15, B => 
                           lpf_filter_inst_lpf_q_n144, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_n167);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_16 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_16, B => 
                           lpf_filter_inst_lpf_q_n143, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_n166);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_17 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_17, B => 
                           lpf_filter_inst_lpf_q_n142, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_n165);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_18 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_18, B => 
                           lpf_filter_inst_lpf_q_n141, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_q_n164);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_19 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_19, B => 
                           lpf_filter_inst_lpf_q_n140, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_q_n163);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_20 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_20, B => 
                           lpf_filter_inst_lpf_q_n139, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_q_n162);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_21 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_21, B => 
                           lpf_filter_inst_lpf_q_n138, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_q_n161);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_22 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_22, B => 
                           lpf_filter_inst_lpf_q_n137, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_23_port, S 
                           => lpf_filter_inst_lpf_q_n160);
   lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_U1_23 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_t12_13_22, B => 
                           lpf_filter_inst_lpf_q_n137, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_carry_23_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_0_root_add_292_n_1104, S 
                           => lpf_filter_inst_lpf_q_n159);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U17 : EXOR2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n15, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n16, Z 
                           => lpf_filter_inst_lpf_q_n92);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U16 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_2, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n14);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U15 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_1, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n15);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U14 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_3, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n13);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U13 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_n117, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n16);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U12 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_14, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U11 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_13, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n3);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U10 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_12, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n4);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U9 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_11, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n5);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U8 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_10, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n6);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U7 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_9, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n7);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U6 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_8, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n8);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U5 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_7, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n9);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U4 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_6, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n10);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U3 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_5, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n11);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_t0_1_4, Z => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n12);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U1 : AND2D1 port map( A1
                           => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n15, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n16, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n1);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_2 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n136, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n14, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n1, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_n91);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_3 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n135, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n13, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_n90);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_4 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n134, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n12, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_n89);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_5 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n133, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n11, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_n88);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_6 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n132, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n10, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_n87);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_7 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n131, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n9, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_n86);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_8 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n130, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n8, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_n85);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_9 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n129, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n7, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_n84);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_10 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n128, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n6, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_n83);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_11 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n127, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n5, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_n194);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_12 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n126, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n4, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_n193);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_13 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n125, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n3, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_n192);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_14 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n124, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_n191);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_15 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n123, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_n190);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_16 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n122, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_n189);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_17 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n121, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_n188);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_18 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n120, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_q_n187);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_19 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n119, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_q_n186);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_20 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n118, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_q_n185);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_21 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n118, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_q_n184);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_22 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n118, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_23_port, S 
                           => lpf_filter_inst_lpf_q_n183);
   lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_U2_23 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n118, B => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n2, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_carry_23_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_3_root_sub_0_root_add_292_n_1109, S 
                           => lpf_filter_inst_lpf_q_n182);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U2 : EXOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_q_n181, A2 => 
                           lpf_filter_inst_lpf_q_n92, Z => 
                           lpf_filter_inst_lpf_q_n116);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1 : AND2D1 port map( A1
                           => lpf_filter_inst_lpf_q_n181, A2 => 
                           lpf_filter_inst_lpf_q_n92, Z => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_n1);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_2 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n91, B => 
                           lpf_filter_inst_lpf_q_n180, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_n1, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_n115);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_3 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n90, B => 
                           lpf_filter_inst_lpf_q_n179, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_n114);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_4 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n89, B => 
                           lpf_filter_inst_lpf_q_n178, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_n113);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_5 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n88, B => 
                           lpf_filter_inst_lpf_q_n177, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_n112);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_6 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n87, B => 
                           lpf_filter_inst_lpf_q_n176, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_n111);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_7 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n86, B => 
                           lpf_filter_inst_lpf_q_n175, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_n110);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_8 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n85, B => 
                           lpf_filter_inst_lpf_q_n174, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_n109);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_9 : ADFULD1 port map(
                           A => lpf_filter_inst_lpf_q_n84, B => 
                           lpf_filter_inst_lpf_q_n173, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_n108);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_10 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n83, B => 
                           lpf_filter_inst_lpf_q_n172, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_n107);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_11 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n194, B => 
                           lpf_filter_inst_lpf_q_n171, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_n106);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_12 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n193, B => 
                           lpf_filter_inst_lpf_q_n170, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_n105);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_13 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n192, B => 
                           lpf_filter_inst_lpf_q_n169, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_n104);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_14 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n191, B => 
                           lpf_filter_inst_lpf_q_n168, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_n103);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_15 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n190, B => 
                           lpf_filter_inst_lpf_q_n167, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_n102);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_16 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n189, B => 
                           lpf_filter_inst_lpf_q_n166, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_n101);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_17 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n188, B => 
                           lpf_filter_inst_lpf_q_n165, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_n100);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_18 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n187, B => 
                           lpf_filter_inst_lpf_q_n164, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_19_port, S 
                           => lpf_filter_inst_lpf_q_n99);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_19 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n186, B => 
                           lpf_filter_inst_lpf_q_n163, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_20_port, S 
                           => lpf_filter_inst_lpf_q_n98);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_20 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n185, B => 
                           lpf_filter_inst_lpf_q_n162, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_21_port, S 
                           => lpf_filter_inst_lpf_q_n97);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_21 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n184, B => 
                           lpf_filter_inst_lpf_q_n161, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_22_port, S 
                           => lpf_filter_inst_lpf_q_n96);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_22 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n183, B => 
                           lpf_filter_inst_lpf_q_n160, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_23_port, S 
                           => lpf_filter_inst_lpf_q_n95);
   lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_U1_23 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n182, B => 
                           lpf_filter_inst_lpf_q_n159, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_carry_23_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_0_root_add_292_n_1113, S 
                           => lpf_filter_inst_lpf_q_n94);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U30 : NOR2M1D1 port map(
                           A1 => lpf_filter_inst_lpf_q_pair0_28_0, A2 => 
                           lpf_filter_inst_lpf_q_n117, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n28);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U29 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n28, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n7, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n29);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U28 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n28, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n7, 
                           B1 => lpf_filter_inst_lpf_q_pair0_28_1, B2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n29, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n26);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U27 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_q_n115, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n26, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n27);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U26 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n26, 
                           B2 => lpf_filter_inst_lpf_q_n115, A1 => 
                           lpf_filter_inst_lpf_q_pair0_28_2, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n27, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n24);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U25 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n24, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n6, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n25);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U24 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n24, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n6, 
                           B1 => lpf_filter_inst_lpf_q_pair0_28_3, B2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n25, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n22);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U23 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_q_n113, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n22, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n23);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U22 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n22, 
                           B2 => lpf_filter_inst_lpf_q_n113, A1 => 
                           lpf_filter_inst_lpf_q_pair0_28_4, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n23, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n20);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U21 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n20, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n5, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n21);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U20 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n20, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n5, 
                           B1 => lpf_filter_inst_lpf_q_pair0_28_5, B2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n21, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n18);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U19 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_q_n111, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n18, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n19);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U18 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n18, 
                           B2 => lpf_filter_inst_lpf_q_n111, A1 => 
                           lpf_filter_inst_lpf_q_pair0_28_6, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n19, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n16);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U17 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n16, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n4, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n17);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U16 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n16, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n4, 
                           B1 => lpf_filter_inst_lpf_q_pair0_28_7, B2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n17, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n14);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U15 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_q_n109, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n14, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n15);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U14 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n14, 
                           B2 => lpf_filter_inst_lpf_q_n109, A1 => 
                           lpf_filter_inst_lpf_q_pair0_28_8, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n15, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n12);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U13 : AND2D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n12, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n3, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n13);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U12 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n12, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n3, 
                           B1 => lpf_filter_inst_lpf_q_pair0_28_9, B2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n13, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n10);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U11 : NOR2D1 port map( 
                           A1 => lpf_filter_inst_lpf_q_n107, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n10, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n11);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U10 : AOI22M20D1 port 
                           map( B1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n10, 
                           B2 => lpf_filter_inst_lpf_q_n107, A1 => 
                           lpf_filter_inst_lpf_q_pair0_28_10, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n11, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n8);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U9 : AND2D1 port map( A1
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n8, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n2, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n9);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U8 : OAI22D1 port map( 
                           A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n8, 
                           A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n2, 
                           B1 => lpf_filter_inst_lpf_q_pair0_28_11, B2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n9, Z 
                           => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_12_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U7 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_pair0_28_12, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U6 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_n108, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n3);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U5 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_n110, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n4);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U4 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_n112, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n5);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U3 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_n114, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n6);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_n116, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n7);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U1 : INVD1 port map( A 
                           => lpf_filter_inst_lpf_q_n106, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n2);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_12 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n105, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_13_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_12_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_13 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n104, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_14_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_13_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_14 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n103, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_15_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_14_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_15 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n102, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_16_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_15_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_16 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n101, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_17_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_16_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_17 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n100, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_18_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_17_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_18 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n99, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_19_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_18_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_19 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n98, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_20_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_19_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_20 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n97, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_20_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_21_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_20_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_21 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n96, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_21_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_22_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_21_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_22 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n95, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_22_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_23_port, S 
                           => 
                           lpf_filter_inst_lpf_q_t0_1_3_4_5_7_8_9_11_12_13_14_22_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_U2_23 : ADFULD1 port 
                           map( A => lpf_filter_inst_lpf_q_n94, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n1, 
                           CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_carry_23_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_0_root_add_292_n_1128, S 
                           => filter_out_q_4_port);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_p206_2_3_port, A2 => 
                           lpf_filter_inst_lpf_q_p206_1_3, Z => 
                           lpf_filter_inst_lpf_q_p206_1_6);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_p206_2_3_port, A2 => 
                           lpf_filter_inst_lpf_q_p206_1_3, Z => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_n1);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_1_4, B => 
                           lpf_filter_inst_lpf_q_p206_2_4_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_n1, CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_7);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_2_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_5_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_8);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_3_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_6_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_9);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_4_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_7_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_10);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_5_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_8_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_11);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_6_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_9_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_12);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_7_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_10_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_13);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_8_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_11_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_14);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_9_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_12_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_15);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_10_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_13_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_16);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair13_15_11_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_14_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_17);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_2_15_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_15_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_19_port, S 
                           => lpf_filter_inst_lpf_q_p206_1_18);
   lpf_filter_inst_lpf_q_add_1_root_add_285_U1_19 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_p206_2_15_port, B => 
                           lpf_filter_inst_lpf_q_p206_2_15_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_carry_19_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_285_n_1158, S 
                           => lpf_filter_inst_lpf_q_p206_1_19);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_60_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_275_port, Z => 
                           lpf_filter_inst_lpf_q_pair4_24_0);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_60_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_275_port, Z => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_n1);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_276_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_61_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_n1, CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_2_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_1);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_277_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_62_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_2);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_278_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_63_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_3);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_279_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_64_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_4);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_280_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_65_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_5);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_281_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_66_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_6);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_282_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_67_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_7);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_283_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_68_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_8);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_284_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_69_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_9);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_285_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_70_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_10);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_286_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_71_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_pair4_24_11);
   lpf_filter_inst_lpf_q_add_2_root_sub_287_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_286_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_71_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_sub_287_n_1268, S 
                           => lpf_filter_inst_lpf_q_pair4_24_12);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_48_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_287_port, Z => 
                           lpf_filter_inst_lpf_q_pair5_23_0);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_48_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_287_port, Z => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_n1);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_288_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_49_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_n1, CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_2_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_1);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_289_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_50_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_2);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_290_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_51_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_3);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_291_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_52_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_4);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_292_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_53_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_5);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_293_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_54_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_6);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_294_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_55_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_7);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_295_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_56_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_8);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_296_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_57_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_9);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_297_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_58_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_10);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_298_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_59_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_pair5_23_11);
   lpf_filter_inst_lpf_q_add_3_root_sub_287_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_298_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_59_port, CI => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_3_root_sub_287_n_1271, S 
                           => lpf_filter_inst_lpf_q_pair5_23_12);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair4_24_0, A2 => 
                           lpf_filter_inst_lpf_q_pair5_23_0, Z => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_3_port);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair4_24_0, A2 => 
                           lpf_filter_inst_lpf_q_pair5_23_0, Z => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_n1);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_1, B => 
                           lpf_filter_inst_lpf_q_pair4_24_1, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_n1, CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_2_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_4_port);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_2, B => 
                           lpf_filter_inst_lpf_q_pair4_24_2, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_2);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_3, B => 
                           lpf_filter_inst_lpf_q_pair4_24_3, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_3);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_4, B => 
                           lpf_filter_inst_lpf_q_pair4_24_4, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_4);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_5, B => 
                           lpf_filter_inst_lpf_q_pair4_24_5, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_5);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_6, B => 
                           lpf_filter_inst_lpf_q_pair4_24_6, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_6);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_7, B => 
                           lpf_filter_inst_lpf_q_pair4_24_7, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_7);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_8, B => 
                           lpf_filter_inst_lpf_q_pair4_24_8, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_9, B => 
                           lpf_filter_inst_lpf_q_pair4_24_9, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_9);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_10, B => 
                           lpf_filter_inst_lpf_q_pair4_24_10, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_10);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_11, B => 
                           lpf_filter_inst_lpf_q_pair4_24_11, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_11);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_12, B => 
                           lpf_filter_inst_lpf_q_pair4_24_12, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_12);
   lpf_filter_inst_lpf_q_add_1_root_sub_287_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair5_23_12, B => 
                           lpf_filter_inst_lpf_q_pair4_24_12, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_287_n_1274, S 
                           => lpf_filter_inst_lpf_q_t4_5_13);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U17 : EXNOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n15, A2 => 
                           lpf_filter_inst_lpf_q_t4_5_2, Z => 
                           lpf_filter_inst_lpf_q_t4_5_8_9_5_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U16 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_0_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n15);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U15 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_13_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n2);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U14 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_2, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n1);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U13 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_10_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n5);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U12 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_9_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n6);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U11 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_8_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n7);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U10 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_7_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n8);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U9 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_6_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n9);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U8 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_5_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n10);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U7 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_4_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n11);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U6 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_3_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n12);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U5 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_2_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n13);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U4 : NAN2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t8_9_0_port, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n1, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_3_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U3 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_1_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n14);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_12_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n3);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U1 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t8_9_11_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n4);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_3, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n14, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_6_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_4, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n13, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_7_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_5, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n12, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_8_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_6, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n11, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_9_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_7, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n10, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_10_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_8, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n9, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_11_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_9, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n8, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_12_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_10, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n7, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_13_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_11, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n6, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_14_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_12, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n5, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_15_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_13, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n4, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_16_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_13, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n3, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_17_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_13, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n2, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_18_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_287_U2_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_t4_5_13, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n2, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_287_n_1279, S 
                           => lpf_filter_inst_lpf_q_t4_5_8_9_19_port);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t11_14_0_port, A2 => 
                           lpf_filter_inst_lpf_q_pair11_17_2_port, Z => 
                           lpf_filter_inst_lpf_q_n66);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_t11_14_0_port, A2 => 
                           lpf_filter_inst_lpf_q_pair11_17_2_port, Z => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_n1);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_3_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_168_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_n1, CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_n65);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_4_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_169_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_n64);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_5_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_170_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_n63);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_6_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_171_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_n82);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_7_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_172_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_n81);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_8_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_173_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_n80);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_9_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_174_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_n79);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_10_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_175_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_n78);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_11_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_176_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_n77);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_12_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_177_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_n76);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_12_port, B => 
                           lpf_filter_inst_lpf_q_p232_2_17, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_n75);
   lpf_filter_inst_lpf_q_add_2_root_add_286_U1_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair11_17_12_port, B => 
                           lpf_filter_inst_lpf_q_p232_2_17, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_286_n_1208, S 
                           => lpf_filter_inst_lpf_q_n62);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U22 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n19, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n20, Z => 
                           lpf_filter_inst_lpf_q_t11_14_1_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U21 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n18, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n2, Z => 
                           lpf_filter_inst_lpf_q_t11_14_2_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U20 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_1, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n19);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U19 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_t11_14_0_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n20);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U18 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_5, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n15);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U17 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_3, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n17);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U16 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n19, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n20, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n2);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U15 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_2, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n18);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U14 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_17, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n3);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U13 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_17, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n4);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U12 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_17, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n5);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U11 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_17, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n6);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U10 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_17, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n7);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U9 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_12, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n8);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U8 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_11, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n9);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U7 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_10, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n10);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U6 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_9, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n11);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U5 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_8, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n12);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U4 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_7, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n13);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U3 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_6, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n14);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_p232_2_4, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n16);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n18, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n2, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n1);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n74, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n17, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n1, CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_3_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n67, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n16, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_4_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n66, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n15, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_5_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n65, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n14, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_6_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n64, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n13, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_7_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n63, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n12, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_8_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n82, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n11, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_9_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n81, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n10, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_10_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n80, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n9, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_11_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n79, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n8, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_12_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n78, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n7, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_13_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n77, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n6, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_14_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n76, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n5, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_16_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_15_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_16 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n75, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n4, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_16_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_17_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_16_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_17 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n62, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n3, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_17_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_18_port, S 
                           => lpf_filter_inst_lpf_q_t11_14_17_port);
   lpf_filter_inst_lpf_q_sub_0_root_add_286_U2_18 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_n62, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n3, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_carry_18_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_add_286_n_1214, S 
                           => lpf_filter_inst_lpf_q_t11_14_18_port);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_108_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_227_port, Z => 
                           lpf_filter_inst_lpf_q_pair8_20_0);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_108_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_227_port, Z => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_n1);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_228_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_109_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_n1, CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_2_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_1);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_229_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_110_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_2);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_230_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_111_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_3);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_231_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_112_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_4);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_232_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_113_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_5);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_233_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_114_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_6);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_234_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_115_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_7);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_235_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_116_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_8);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_236_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_117_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_9);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_237_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_118_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_10);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_238_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_119_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_pair8_20_11);
   lpf_filter_inst_lpf_q_add_1_root_add_277_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_238_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_119_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_add_277_n_1290, S 
                           => lpf_filter_inst_lpf_q_pair8_20_12);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_96_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_239_port, Z => 
                           lpf_filter_inst_lpf_q_pair9_19_0);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_96_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_239_port, Z => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_n1);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_240_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_97_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_n1, CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_2_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_1);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_241_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_98_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_2);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_242_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_99_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_3);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_243_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_100_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_4);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_244_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_101_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_5);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_245_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_102_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_6);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_246_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_103_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_7);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_247_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_104_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_8);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_248_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_105_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_9);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_249_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_106_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_10);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_250_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_107_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_pair9_19_11);
   lpf_filter_inst_lpf_q_add_2_root_add_277_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_250_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_107_port, CI => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_2_root_add_277_n_1293, S 
                           => lpf_filter_inst_lpf_q_pair9_19_12);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair8_20_0, A2 => 
                           lpf_filter_inst_lpf_q_pair9_19_0, Z => 
                           lpf_filter_inst_lpf_q_t8_9_0_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair8_20_0, A2 => 
                           lpf_filter_inst_lpf_q_pair9_19_0, Z => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_n1);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_13 : EXOR3D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair9_19_12, A2 => 
                           lpf_filter_inst_lpf_q_pair8_20_12, A3 => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_13_port, Z 
                           => lpf_filter_inst_lpf_q_t8_9_13_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_1, B => 
                           lpf_filter_inst_lpf_q_pair8_20_1, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_n1, CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_2_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_1_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_2, B => 
                           lpf_filter_inst_lpf_q_pair8_20_2, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_2_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_3, B => 
                           lpf_filter_inst_lpf_q_pair8_20_3, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_3_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_4, B => 
                           lpf_filter_inst_lpf_q_pair8_20_4, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_4_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_5, B => 
                           lpf_filter_inst_lpf_q_pair8_20_5, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_5_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_6, B => 
                           lpf_filter_inst_lpf_q_pair8_20_6, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_6_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_7, B => 
                           lpf_filter_inst_lpf_q_pair8_20_7, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_7_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_8, B => 
                           lpf_filter_inst_lpf_q_pair8_20_8, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_8_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_9, B => 
                           lpf_filter_inst_lpf_q_pair8_20_9, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_9_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_10, B => 
                           lpf_filter_inst_lpf_q_pair8_20_10, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_10_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_11, B => 
                           lpf_filter_inst_lpf_q_pair8_20_11, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_11_port);
   lpf_filter_inst_lpf_q_add_0_root_add_277_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair9_19_12, B => 
                           lpf_filter_inst_lpf_q_pair8_20_12, CI => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_0_root_add_277_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_t8_9_12_port);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U2 : EXOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_36_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_299_port, Z => 
                           lpf_filter_inst_lpf_q_n136);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1 : AND2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_36_port, A2 => 
                           lpf_filter_inst_lpf_q_arx_input_reg_299_port, Z => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_n1);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_1 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_300_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_37_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_n1, CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_2_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_1_port);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_2 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_301_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_38_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_2_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_3_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_2);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_302_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_39_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_3);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_303_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_40_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_4);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_304_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_41_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_5);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_305_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_42_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_6);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_306_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_43_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_7);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_307_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_44_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_8);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_308_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_45_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_9);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_309_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_46_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_10);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_310_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_47_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_pair3_25_11);
   lpf_filter_inst_lpf_q_add_1_root_sub_279_U1_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_arx_input_reg_310_port, B => 
                           lpf_filter_inst_lpf_q_arx_input_reg_47_port, CI => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_add_1_root_sub_279_n_1189, S 
                           => lpf_filter_inst_lpf_q_pair3_25_12);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U16 : EXNOR2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n14, A2 => 
                           lpf_filter_inst_lpf_q_pair3_25_2, Z => 
                           lpf_filter_inst_lpf_q_t3_7_2_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U15 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_0_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n14);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U14 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_12_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n2);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U13 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_2, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n1);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U12 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_9_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n5);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U11 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_8_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n6);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U10 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_7_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n7);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U9 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_6_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n8);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U8 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_5_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n9);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U7 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_4_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n10);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U6 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_3_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n11);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U5 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_2_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n12);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U4 : NAN2D1 port map( A1 => 
                           lpf_filter_inst_lpf_q_pair7_21_0_port, A2 => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n1, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_3_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U3 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_1_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n13);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_11_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n3);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U1 : INVD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair7_21_10_port, Z => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n4);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_3 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_3, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n13, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_3_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_4_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_3_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_4 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_4, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n12, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_4_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_5_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_4_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_5 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_5, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n11, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_5_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_6_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_5_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_6 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_6, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n10, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_6_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_7_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_6_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_7 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_7, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n9, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_7_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_8_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_7_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_8 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_8, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n8, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_8_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_9_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_8_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_9 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_9, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n7, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_9_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_10_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_9_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_10 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_10, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n6, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_10_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_11_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_10_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_11 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_11, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n5, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_11_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_12_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_11_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_12 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_12, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n4, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_12_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_13_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_12_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_13 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_12, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n3, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_13_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_14_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_13_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_14 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_12, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n2, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_14_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_15_port, S 
                           => lpf_filter_inst_lpf_q_t3_7_14_port);
   lpf_filter_inst_lpf_q_sub_0_root_sub_279_U2_15 : ADFULD1 port map( A => 
                           lpf_filter_inst_lpf_q_pair3_25_12, B => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n2, CI => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_carry_15_port, 
                           CO => 
                           lpf_filter_inst_lpf_q_sub_0_root_sub_279_n_1194, S 
                           => lpf_filter_inst_lpf_q_t3_7_15_port);
   dam_demodulator_inst_U18 : TIELO port map( Z => dam_demodulator_inst_n10);
   dam_demodulator_inst_U17 : INVD1 port map( A => clk4, Z => 
                           dam_demodulator_inst_n6);
   dam_demodulator_inst_U16 : INVD1 port map( A => rstn, Z => 
                           dam_demodulator_inst_n9);
   dam_demodulator_inst_U15 : OAI21M20D1 port map( A1 => 
                           dam_demodulator_inst_arx_result_reg_2_port, A2 => 
                           dam_demodulator_inst_n2, B => 
                           dam_demodulator_inst_n3, Z => demodulator_out_0_port
                           );
   dam_demodulator_inst_U14 : OAI21M20D1 port map( A1 => 
                           dam_demodulator_inst_arx_result_reg_7_port, A2 => 
                           dam_demodulator_inst_n2, B => 
                           dam_demodulator_inst_n3, Z => demodulator_out_5_port
                           );
   dam_demodulator_inst_U13 : OAI21M20D1 port map( A1 => 
                           dam_demodulator_inst_arx_result_reg_6_port, A2 => 
                           dam_demodulator_inst_n2, B => 
                           dam_demodulator_inst_n3, Z => demodulator_out_4_port
                           );
   dam_demodulator_inst_U12 : OAI21M20D1 port map( A1 => 
                           dam_demodulator_inst_arx_result_reg_5_port, A2 => 
                           dam_demodulator_inst_n2, B => 
                           dam_demodulator_inst_n3, Z => demodulator_out_3_port
                           );
   dam_demodulator_inst_U9 : OAI21M20D1 port map( A1 => 
                           dam_demodulator_inst_arx_result_reg_4_port, A2 => 
                           dam_demodulator_inst_n2, B => 
                           dam_demodulator_inst_n3, Z => demodulator_out_2_port
                           );
   dam_demodulator_inst_U8 : OAI21M20D1 port map( A1 => 
                           dam_demodulator_inst_arx_result_reg_3_port, A2 => 
                           dam_demodulator_inst_n2, B => 
                           dam_demodulator_inst_n3, Z => demodulator_out_1_port
                           );
   dam_demodulator_inst_U7 : NAN3D1 port map( A1 => 
                           dam_demodulator_inst_arx_result_reg_8_port, A2 => 
                           demodulator_out_6_port, A3 => 
                           dam_demodulator_inst_arx_result_reg_9_port, Z => 
                           dam_demodulator_inst_n4);
   dam_demodulator_inst_U6 : INVD1 port map( A => dam_demodulator_inst_n6, Z =>
                           dam_demodulator_inst_n5);
   dam_demodulator_inst_U5 : INVD1 port map( A => dam_demodulator_inst_n6, Z =>
                           dam_demodulator_inst_n1);
   dam_demodulator_inst_U4 : INVD1 port map( A => dam_demodulator_inst_n9, Z =>
                           dam_demodulator_inst_n8);
   dam_demodulator_inst_U3 : INVD1 port map( A => dam_demodulator_inst_n9, Z =>
                           dam_demodulator_inst_n7);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_1_3 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_18_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_13_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_1_4 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_19_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_14_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_0_0 : DFFRPQ1 port map( D => 
                           filter_out_q_0_port, CK => dam_demodulator_inst_n1, 
                           RB => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_15_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_0_1 : DFFRPQ1 port map( D => 
                           filter_out_q_1_port, CK => dam_demodulator_inst_n5, 
                           RB => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_16_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_0_2 : DFFRPQ1 port map( D => 
                           filter_out_q_2_port, CK => dam_demodulator_inst_n1, 
                           RB => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_17_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_0_3 : DFFRPQ1 port map( D => 
                           filter_out_q_3_port, CK => dam_demodulator_inst_n5, 
                           RB => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_18_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_0_4 : DFFRPQ1 port map( D => 
                           filter_out_q_4_port, CK => dam_demodulator_inst_n1, 
                           RB => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_19_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_2_0 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_10_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_5_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_2_1 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_11_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_6_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_2_2 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_12_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_7_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_2_3 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_13_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_8_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_2_4 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_14_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_9_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_1_0 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_15_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_10_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_1_1 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_16_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_11_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_1_2 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_17_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_12_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_1_3 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_18_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_13_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_1_4 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_19_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_14_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_0_0 : DFFRPQ1 port map( D => 
                           filter_out_i_0_port, CK => dam_demodulator_inst_n5, 
                           RB => dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_15_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_0_1 : DFFRPQ1 port map( D => 
                           filter_out_i_1_port, CK => clk4, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_16_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_0_2 : DFFRPQ1 port map( D => 
                           filter_out_i_2_port, CK => clk4, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_17_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_0_3 : DFFRPQ1 port map( D => 
                           filter_out_i_3_port, CK => clk4, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_18_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_0_4 : DFFRPQ1 port map( D => 
                           filter_out_i_4_port, CK => clk4, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_19_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_2_0 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_10_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_5_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_2_1 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_11_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_6_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_2_2 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_12_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_7_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_2_3 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_13_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_8_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_2_4 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_14_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_9_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_1_0 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_15_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_10_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_1_1 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_16_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_11_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_1_2 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_17_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_12_port);
   dam_demodulator_inst_arx_result_reg_reg_10 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_10_port, CK => clk4, RB 
                           => dam_demodulator_inst_n8, Q => 
                           demodulator_out_6_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_3_4 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_9_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_4_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_3_4 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_9_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_4_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_3_2 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_7_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_2_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_3_3 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_8_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_3_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_3_2 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_7_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_2_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_3_3 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_8_port, 
                           CK => dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_3_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_3_0 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_5_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_0_port);
   dam_demodulator_inst_arx_dem_samples_q_reg_reg_3_1 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_6_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_1_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_3_0 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_5_port, 
                           CK => dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_0_port);
   dam_demodulator_inst_arx_dem_samples_i_reg_reg_3_1 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_6_port, 
                           CK => clk4, RB => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_1_port);
   dam_demodulator_inst_arx_result_reg_reg_9 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_9_port, CK => clk4, RB 
                           => dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_result_reg_9_port);
   dam_demodulator_inst_arx_result_reg_reg_8 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_8_port, CK => clk4, RB 
                           => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_result_reg_8_port);
   dam_demodulator_inst_arx_result_reg_reg_2 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_2_port, CK => clk4, RB 
                           => dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_result_reg_2_port);
   dam_demodulator_inst_arx_result_reg_reg_3 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_3_port, CK => clk4, RB 
                           => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_result_reg_3_port);
   dam_demodulator_inst_arx_result_reg_reg_4 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_4_port, CK => clk4, RB 
                           => dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_result_reg_4_port);
   dam_demodulator_inst_arx_result_reg_reg_5 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_5_port, CK => 
                           dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_result_reg_5_port);
   dam_demodulator_inst_arx_result_reg_reg_6 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_6_port, CK => 
                           dam_demodulator_inst_n1, RB => 
                           dam_demodulator_inst_n8, Q => 
                           dam_demodulator_inst_arx_result_reg_6_port);
   dam_demodulator_inst_arx_result_reg_reg_7 : DFFRPQ1 port map( D => 
                           dam_demodulator_inst_result_7_port, CK => 
                           dam_demodulator_inst_n5, RB => 
                           dam_demodulator_inst_n7, Q => 
                           dam_demodulator_inst_arx_result_reg_7_port);
   dam_demodulator_inst_U11 : OAI31D1 port map( A1 => demodulator_out_6_port, 
                           A2 => dam_demodulator_inst_arx_result_reg_9_port, A3
                           => dam_demodulator_inst_arx_result_reg_8_port, B => 
                           dam_demodulator_inst_n4, Z => 
                           dam_demodulator_inst_n2);
   dam_demodulator_inst_U10 : OR2D1 port map( A1 => dam_demodulator_inst_n2, A2
                           => demodulator_out_6_port, Z => 
                           dam_demodulator_inst_n3);
   dam_demodulator_inst_mult_131_U95 : NAN2D1 port map( A1 => 
                           filter_out_i_2_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_3_port, Z
                           => dam_demodulator_inst_mult_131_n101);
   dam_demodulator_inst_mult_131_U94 : NAN2D1 port map( A1 => 
                           filter_out_i_3_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_2_port, Z
                           => dam_demodulator_inst_mult_131_n100);
   dam_demodulator_inst_mult_131_U93 : NAN2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n101, A2 => 
                           dam_demodulator_inst_mult_131_n100, Z => 
                           dam_demodulator_inst_mult_131_n19);
   dam_demodulator_inst_mult_131_U92 : EXNOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n100, A2 => 
                           dam_demodulator_inst_mult_131_n101, Z => 
                           dam_demodulator_inst_mult_131_n20);
   dam_demodulator_inst_mult_131_U91 : AND2D1 port map( A1 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_4_port, 
                           A2 => filter_out_i_4_port, Z => 
                           dam_demodulator_inst_mult_131_n33);
   dam_demodulator_inst_mult_131_U90 : NAN2D1 port map( A1 => 
                           filter_out_i_4_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_3_port, Z
                           => dam_demodulator_inst_mult_131_n34);
   dam_demodulator_inst_mult_131_U89 : NAN2D1 port map( A1 => 
                           filter_out_i_4_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_2_port, Z
                           => dam_demodulator_inst_mult_131_n35);
   dam_demodulator_inst_mult_131_U88 : NAN2D1 port map( A1 => 
                           filter_out_i_4_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_1_port, Z
                           => dam_demodulator_inst_mult_131_n36);
   dam_demodulator_inst_mult_131_U87 : NAN2D1 port map( A1 => 
                           filter_out_i_4_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_0_port, Z
                           => dam_demodulator_inst_mult_131_n37);
   dam_demodulator_inst_mult_131_U86 : NAN2D1 port map( A1 => 
                           filter_out_i_3_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_4_port, Z
                           => dam_demodulator_inst_mult_131_n38);
   dam_demodulator_inst_mult_131_U85 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n96, A2 => 
                           dam_demodulator_inst_mult_131_n95, Z => 
                           dam_demodulator_inst_mult_131_n39);
   dam_demodulator_inst_mult_131_U84 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n98, A2 => 
                           dam_demodulator_inst_mult_131_n95, Z => 
                           dam_demodulator_inst_mult_131_n41);
   dam_demodulator_inst_mult_131_U83 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n99, A2 => 
                           dam_demodulator_inst_mult_131_n95, Z => 
                           dam_demodulator_inst_mult_131_n42);
   dam_demodulator_inst_mult_131_U82 : NAN2D1 port map( A1 => 
                           filter_out_i_2_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_4_port, Z
                           => dam_demodulator_inst_mult_131_n43);
   dam_demodulator_inst_mult_131_U81 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n97, A2 => 
                           dam_demodulator_inst_mult_131_n94, Z => 
                           dam_demodulator_inst_mult_131_n45);
   dam_demodulator_inst_mult_131_U80 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n98, A2 => 
                           dam_demodulator_inst_mult_131_n94, Z => 
                           dam_demodulator_inst_mult_131_n46);
   dam_demodulator_inst_mult_131_U79 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n99, A2 => 
                           dam_demodulator_inst_mult_131_n94, Z => 
                           dam_demodulator_inst_mult_131_n47);
   dam_demodulator_inst_mult_131_U78 : NAN2D1 port map( A1 => 
                           filter_out_i_1_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_4_port, Z
                           => dam_demodulator_inst_mult_131_n48);
   dam_demodulator_inst_mult_131_U77 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n96, A2 => 
                           dam_demodulator_inst_mult_131_n93, Z => 
                           dam_demodulator_inst_mult_131_n49);
   dam_demodulator_inst_mult_131_U76 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n97, A2 => 
                           dam_demodulator_inst_mult_131_n93, Z => 
                           dam_demodulator_inst_mult_131_n50);
   dam_demodulator_inst_mult_131_U75 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n98, A2 => 
                           dam_demodulator_inst_mult_131_n93, Z => 
                           dam_demodulator_inst_mult_131_n51);
   dam_demodulator_inst_mult_131_U74 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n99, A2 => 
                           dam_demodulator_inst_mult_131_n93, Z => 
                           dam_demodulator_inst_mult_131_n52);
   dam_demodulator_inst_mult_131_U73 : NAN2D1 port map( A1 => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_4_port, 
                           A2 => filter_out_i_0_port, Z => 
                           dam_demodulator_inst_mult_131_n53);
   dam_demodulator_inst_mult_131_U72 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n92, A2 => 
                           dam_demodulator_inst_mult_131_n96, Z => 
                           dam_demodulator_inst_mult_131_n54);
   dam_demodulator_inst_mult_131_U71 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n92, A2 => 
                           dam_demodulator_inst_mult_131_n97, Z => 
                           dam_demodulator_inst_mult_131_n55);
   dam_demodulator_inst_mult_131_U70 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n92, A2 => 
                           dam_demodulator_inst_mult_131_n98, Z => 
                           dam_demodulator_inst_mult_131_n56);
   dam_demodulator_inst_mult_131_U69 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_131_n92, A2 => 
                           dam_demodulator_inst_mult_131_n99, Z => 
                           dam_demodulator_inst_prod_i_qd_0);
   dam_demodulator_inst_mult_131_U68 : INVD1 port map( A => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_3_port, Z
                           => dam_demodulator_inst_mult_131_n96);
   dam_demodulator_inst_mult_131_U67 : INVD1 port map( A => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_2_port, Z
                           => dam_demodulator_inst_mult_131_n97);
   dam_demodulator_inst_mult_131_U66 : INVD1 port map( A => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_0_port, Z
                           => dam_demodulator_inst_mult_131_n99);
   dam_demodulator_inst_mult_131_U65 : INVD1 port map( A => 
                           dam_demodulator_inst_arx_dem_samples_q_reg_1_port, Z
                           => dam_demodulator_inst_mult_131_n98);
   dam_demodulator_inst_mult_131_U64 : INVD1 port map( A => 
                           dam_demodulator_inst_mult_131_n1, Z => 
                           dam_demodulator_inst_prod_i_qd_9);
   dam_demodulator_inst_mult_131_U63 : INVD1 port map( A => filter_out_i_3_port
                           , Z => dam_demodulator_inst_mult_131_n95);
   dam_demodulator_inst_mult_131_U62 : INVD1 port map( A => filter_out_i_2_port
                           , Z => dam_demodulator_inst_mult_131_n94);
   dam_demodulator_inst_mult_131_U61 : INVD1 port map( A => filter_out_i_1_port
                           , Z => dam_demodulator_inst_mult_131_n93);
   dam_demodulator_inst_mult_131_U60 : INVD1 port map( A => filter_out_i_0_port
                           , Z => dam_demodulator_inst_mult_131_n92);
   dam_demodulator_inst_mult_131_U22 : ADHALFDL port map( A => 
                           dam_demodulator_inst_mult_131_n51, B => 
                           dam_demodulator_inst_mult_131_n55, CO => 
                           dam_demodulator_inst_mult_131_n31, S => 
                           dam_demodulator_inst_mult_131_n32);
   dam_demodulator_inst_mult_131_U21 : ADHALFDL port map( A => 
                           dam_demodulator_inst_mult_131_n42, B => 
                           dam_demodulator_inst_mult_131_n46, CO => 
                           dam_demodulator_inst_mult_131_n29, S => 
                           dam_demodulator_inst_mult_131_n30);
   dam_demodulator_inst_mult_131_U20 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n50, B => 
                           dam_demodulator_inst_mult_131_n54, CI => 
                           dam_demodulator_inst_mult_131_n31, CO => 
                           dam_demodulator_inst_mult_131_n27, S => 
                           dam_demodulator_inst_mult_131_n28);
   dam_demodulator_inst_mult_131_U19 : ADHALFDL port map( A => 
                           dam_demodulator_inst_mult_131_n49, B => 
                           dam_demodulator_inst_mult_131_n41, CO => 
                           dam_demodulator_inst_mult_131_n25, S => 
                           dam_demodulator_inst_mult_131_n26);
   dam_demodulator_inst_mult_131_U18 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n53, B => 
                           dam_demodulator_inst_mult_131_n45, CI => 
                           dam_demodulator_inst_mult_131_n37, CO => 
                           dam_demodulator_inst_mult_131_n23, S => 
                           dam_demodulator_inst_mult_131_n24);
   dam_demodulator_inst_mult_131_U17 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n26, B => 
                           dam_demodulator_inst_mult_131_n29, CI => 
                           dam_demodulator_inst_mult_131_n27, CO => 
                           dam_demodulator_inst_mult_131_n21, S => 
                           dam_demodulator_inst_mult_131_n22);
   dam_demodulator_inst_mult_131_U14 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n36, B => 
                           dam_demodulator_inst_mult_131_n48, CI => 
                           dam_demodulator_inst_mult_131_n25, CO => 
                           dam_demodulator_inst_mult_131_n17, S => 
                           dam_demodulator_inst_mult_131_n18);
   dam_demodulator_inst_mult_131_U13 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n23, B => 
                           dam_demodulator_inst_mult_131_n20, CI => 
                           dam_demodulator_inst_mult_131_n18, CO => 
                           dam_demodulator_inst_mult_131_n15, S => 
                           dam_demodulator_inst_mult_131_n16);
   dam_demodulator_inst_mult_131_U12 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n43, B => 
                           dam_demodulator_inst_mult_131_n39, CI => 
                           dam_demodulator_inst_mult_131_n35, CO => 
                           dam_demodulator_inst_mult_131_n13, S => 
                           dam_demodulator_inst_mult_131_n14);
   dam_demodulator_inst_mult_131_U11 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n17, B => 
                           dam_demodulator_inst_mult_131_n19, CI => 
                           dam_demodulator_inst_mult_131_n14, CO => 
                           dam_demodulator_inst_mult_131_n11, S => 
                           dam_demodulator_inst_mult_131_n12);
   dam_demodulator_inst_mult_131_U10 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n34, B => 
                           dam_demodulator_inst_mult_131_n38, CI => 
                           dam_demodulator_inst_mult_131_n13, CO => 
                           dam_demodulator_inst_mult_131_n9, S => 
                           dam_demodulator_inst_mult_131_n10);
   dam_demodulator_inst_mult_131_U9 : ADHALFDL port map( A => 
                           dam_demodulator_inst_mult_131_n56, B => 
                           dam_demodulator_inst_mult_131_n52, CO => 
                           dam_demodulator_inst_mult_131_n8, S => 
                           dam_demodulator_inst_prod_i_qd_1);
   dam_demodulator_inst_mult_131_U8 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n8, B => 
                           dam_demodulator_inst_mult_131_n47, CI => 
                           dam_demodulator_inst_mult_131_n32, CO => 
                           dam_demodulator_inst_mult_131_n7, S => 
                           dam_demodulator_inst_prod_i_qd_2);
   dam_demodulator_inst_mult_131_U7 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n7, B => 
                           dam_demodulator_inst_mult_131_n30, CI => 
                           dam_demodulator_inst_mult_131_n28, CO => 
                           dam_demodulator_inst_mult_131_n6, S => 
                           dam_demodulator_inst_prod_i_qd_3);
   dam_demodulator_inst_mult_131_U6 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n22, B => 
                           dam_demodulator_inst_mult_131_n24, CI => 
                           dam_demodulator_inst_mult_131_n6, CO => 
                           dam_demodulator_inst_mult_131_n5, S => 
                           dam_demodulator_inst_prod_i_qd_4);
   dam_demodulator_inst_mult_131_U5 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n16, B => 
                           dam_demodulator_inst_mult_131_n21, CI => 
                           dam_demodulator_inst_mult_131_n5, CO => 
                           dam_demodulator_inst_mult_131_n4, S => 
                           dam_demodulator_inst_prod_i_qd_5);
   dam_demodulator_inst_mult_131_U4 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n12, B => 
                           dam_demodulator_inst_mult_131_n15, CI => 
                           dam_demodulator_inst_mult_131_n4, CO => 
                           dam_demodulator_inst_mult_131_n3, S => 
                           dam_demodulator_inst_prod_i_qd_6);
   dam_demodulator_inst_mult_131_U3 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n11, B => 
                           dam_demodulator_inst_mult_131_n10, CI => 
                           dam_demodulator_inst_mult_131_n3, CO => 
                           dam_demodulator_inst_mult_131_n2, S => 
                           dam_demodulator_inst_prod_i_qd_7);
   dam_demodulator_inst_mult_131_U2 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_131_n9, B => 
                           dam_demodulator_inst_mult_131_n33, CI => 
                           dam_demodulator_inst_mult_131_n2, CO => 
                           dam_demodulator_inst_mult_131_n1, S => 
                           dam_demodulator_inst_prod_i_qd_8);
   dam_demodulator_inst_mult_130_U95 : NAN2D1 port map( A1 => 
                           filter_out_q_2_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_3_port, Z
                           => dam_demodulator_inst_mult_130_n101);
   dam_demodulator_inst_mult_130_U94 : NAN2D1 port map( A1 => 
                           filter_out_q_3_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_2_port, Z
                           => dam_demodulator_inst_mult_130_n100);
   dam_demodulator_inst_mult_130_U93 : NAN2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n101, A2 => 
                           dam_demodulator_inst_mult_130_n100, Z => 
                           dam_demodulator_inst_mult_130_n19);
   dam_demodulator_inst_mult_130_U92 : EXNOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n100, A2 => 
                           dam_demodulator_inst_mult_130_n101, Z => 
                           dam_demodulator_inst_mult_130_n20);
   dam_demodulator_inst_mult_130_U91 : AND2D1 port map( A1 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_4_port, 
                           A2 => filter_out_q_4_port, Z => 
                           dam_demodulator_inst_mult_130_n33);
   dam_demodulator_inst_mult_130_U90 : NAN2D1 port map( A1 => 
                           filter_out_q_4_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_3_port, Z
                           => dam_demodulator_inst_mult_130_n34);
   dam_demodulator_inst_mult_130_U89 : NAN2D1 port map( A1 => 
                           filter_out_q_4_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_2_port, Z
                           => dam_demodulator_inst_mult_130_n35);
   dam_demodulator_inst_mult_130_U88 : NAN2D1 port map( A1 => 
                           filter_out_q_4_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_1_port, Z
                           => dam_demodulator_inst_mult_130_n36);
   dam_demodulator_inst_mult_130_U87 : NAN2D1 port map( A1 => 
                           filter_out_q_4_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_0_port, Z
                           => dam_demodulator_inst_mult_130_n37);
   dam_demodulator_inst_mult_130_U86 : NAN2D1 port map( A1 => 
                           filter_out_q_3_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_4_port, Z
                           => dam_demodulator_inst_mult_130_n38);
   dam_demodulator_inst_mult_130_U85 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n96, A2 => 
                           dam_demodulator_inst_mult_130_n95, Z => 
                           dam_demodulator_inst_mult_130_n39);
   dam_demodulator_inst_mult_130_U84 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n98, A2 => 
                           dam_demodulator_inst_mult_130_n95, Z => 
                           dam_demodulator_inst_mult_130_n41);
   dam_demodulator_inst_mult_130_U83 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n99, A2 => 
                           dam_demodulator_inst_mult_130_n95, Z => 
                           dam_demodulator_inst_mult_130_n42);
   dam_demodulator_inst_mult_130_U82 : NAN2D1 port map( A1 => 
                           filter_out_q_2_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_4_port, Z
                           => dam_demodulator_inst_mult_130_n43);
   dam_demodulator_inst_mult_130_U81 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n97, A2 => 
                           dam_demodulator_inst_mult_130_n94, Z => 
                           dam_demodulator_inst_mult_130_n45);
   dam_demodulator_inst_mult_130_U80 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n98, A2 => 
                           dam_demodulator_inst_mult_130_n94, Z => 
                           dam_demodulator_inst_mult_130_n46);
   dam_demodulator_inst_mult_130_U79 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n99, A2 => 
                           dam_demodulator_inst_mult_130_n94, Z => 
                           dam_demodulator_inst_mult_130_n47);
   dam_demodulator_inst_mult_130_U78 : NAN2D1 port map( A1 => 
                           filter_out_q_1_port, A2 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_4_port, Z
                           => dam_demodulator_inst_mult_130_n48);
   dam_demodulator_inst_mult_130_U77 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n96, A2 => 
                           dam_demodulator_inst_mult_130_n93, Z => 
                           dam_demodulator_inst_mult_130_n49);
   dam_demodulator_inst_mult_130_U76 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n97, A2 => 
                           dam_demodulator_inst_mult_130_n93, Z => 
                           dam_demodulator_inst_mult_130_n50);
   dam_demodulator_inst_mult_130_U75 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n98, A2 => 
                           dam_demodulator_inst_mult_130_n93, Z => 
                           dam_demodulator_inst_mult_130_n51);
   dam_demodulator_inst_mult_130_U74 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n99, A2 => 
                           dam_demodulator_inst_mult_130_n93, Z => 
                           dam_demodulator_inst_mult_130_n52);
   dam_demodulator_inst_mult_130_U73 : NAN2D1 port map( A1 => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_4_port, 
                           A2 => filter_out_q_0_port, Z => 
                           dam_demodulator_inst_mult_130_n53);
   dam_demodulator_inst_mult_130_U72 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n92, A2 => 
                           dam_demodulator_inst_mult_130_n96, Z => 
                           dam_demodulator_inst_mult_130_n54);
   dam_demodulator_inst_mult_130_U71 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n92, A2 => 
                           dam_demodulator_inst_mult_130_n97, Z => 
                           dam_demodulator_inst_mult_130_n55);
   dam_demodulator_inst_mult_130_U70 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n92, A2 => 
                           dam_demodulator_inst_mult_130_n98, Z => 
                           dam_demodulator_inst_mult_130_n56);
   dam_demodulator_inst_mult_130_U69 : NOR2D1 port map( A1 => 
                           dam_demodulator_inst_mult_130_n92, A2 => 
                           dam_demodulator_inst_mult_130_n99, Z => 
                           dam_demodulator_inst_prod_q_id_0);
   dam_demodulator_inst_mult_130_U68 : INVD1 port map( A => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_3_port, Z
                           => dam_demodulator_inst_mult_130_n96);
   dam_demodulator_inst_mult_130_U67 : INVD1 port map( A => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_2_port, Z
                           => dam_demodulator_inst_mult_130_n97);
   dam_demodulator_inst_mult_130_U66 : INVD1 port map( A => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_0_port, Z
                           => dam_demodulator_inst_mult_130_n99);
   dam_demodulator_inst_mult_130_U65 : INVD1 port map( A => 
                           dam_demodulator_inst_arx_dem_samples_i_reg_1_port, Z
                           => dam_demodulator_inst_mult_130_n98);
   dam_demodulator_inst_mult_130_U64 : INVD1 port map( A => 
                           dam_demodulator_inst_mult_130_n1, Z => 
                           dam_demodulator_inst_prod_q_id_9);
   dam_demodulator_inst_mult_130_U63 : INVD1 port map( A => filter_out_q_3_port
                           , Z => dam_demodulator_inst_mult_130_n95);
   dam_demodulator_inst_mult_130_U62 : INVD1 port map( A => filter_out_q_2_port
                           , Z => dam_demodulator_inst_mult_130_n94);
   dam_demodulator_inst_mult_130_U61 : INVD1 port map( A => filter_out_q_1_port
                           , Z => dam_demodulator_inst_mult_130_n93);
   dam_demodulator_inst_mult_130_U60 : INVD1 port map( A => filter_out_q_0_port
                           , Z => dam_demodulator_inst_mult_130_n92);
   dam_demodulator_inst_mult_130_U22 : ADHALFDL port map( A => 
                           dam_demodulator_inst_mult_130_n51, B => 
                           dam_demodulator_inst_mult_130_n55, CO => 
                           dam_demodulator_inst_mult_130_n31, S => 
                           dam_demodulator_inst_mult_130_n32);
   dam_demodulator_inst_mult_130_U21 : ADHALFDL port map( A => 
                           dam_demodulator_inst_mult_130_n42, B => 
                           dam_demodulator_inst_mult_130_n46, CO => 
                           dam_demodulator_inst_mult_130_n29, S => 
                           dam_demodulator_inst_mult_130_n30);
   dam_demodulator_inst_mult_130_U20 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n50, B => 
                           dam_demodulator_inst_mult_130_n54, CI => 
                           dam_demodulator_inst_mult_130_n31, CO => 
                           dam_demodulator_inst_mult_130_n27, S => 
                           dam_demodulator_inst_mult_130_n28);
   dam_demodulator_inst_mult_130_U19 : ADHALFDL port map( A => 
                           dam_demodulator_inst_mult_130_n49, B => 
                           dam_demodulator_inst_mult_130_n41, CO => 
                           dam_demodulator_inst_mult_130_n25, S => 
                           dam_demodulator_inst_mult_130_n26);
   dam_demodulator_inst_mult_130_U18 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n53, B => 
                           dam_demodulator_inst_mult_130_n45, CI => 
                           dam_demodulator_inst_mult_130_n37, CO => 
                           dam_demodulator_inst_mult_130_n23, S => 
                           dam_demodulator_inst_mult_130_n24);
   dam_demodulator_inst_mult_130_U17 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n26, B => 
                           dam_demodulator_inst_mult_130_n29, CI => 
                           dam_demodulator_inst_mult_130_n27, CO => 
                           dam_demodulator_inst_mult_130_n21, S => 
                           dam_demodulator_inst_mult_130_n22);
   dam_demodulator_inst_mult_130_U14 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n36, B => 
                           dam_demodulator_inst_mult_130_n48, CI => 
                           dam_demodulator_inst_mult_130_n25, CO => 
                           dam_demodulator_inst_mult_130_n17, S => 
                           dam_demodulator_inst_mult_130_n18);
   dam_demodulator_inst_mult_130_U13 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n23, B => 
                           dam_demodulator_inst_mult_130_n20, CI => 
                           dam_demodulator_inst_mult_130_n18, CO => 
                           dam_demodulator_inst_mult_130_n15, S => 
                           dam_demodulator_inst_mult_130_n16);
   dam_demodulator_inst_mult_130_U12 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n43, B => 
                           dam_demodulator_inst_mult_130_n39, CI => 
                           dam_demodulator_inst_mult_130_n35, CO => 
                           dam_demodulator_inst_mult_130_n13, S => 
                           dam_demodulator_inst_mult_130_n14);
   dam_demodulator_inst_mult_130_U11 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n17, B => 
                           dam_demodulator_inst_mult_130_n19, CI => 
                           dam_demodulator_inst_mult_130_n14, CO => 
                           dam_demodulator_inst_mult_130_n11, S => 
                           dam_demodulator_inst_mult_130_n12);
   dam_demodulator_inst_mult_130_U10 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n34, B => 
                           dam_demodulator_inst_mult_130_n38, CI => 
                           dam_demodulator_inst_mult_130_n13, CO => 
                           dam_demodulator_inst_mult_130_n9, S => 
                           dam_demodulator_inst_mult_130_n10);
   dam_demodulator_inst_mult_130_U9 : ADHALFDL port map( A => 
                           dam_demodulator_inst_mult_130_n56, B => 
                           dam_demodulator_inst_mult_130_n52, CO => 
                           dam_demodulator_inst_mult_130_n8, S => 
                           dam_demodulator_inst_prod_q_id_1);
   dam_demodulator_inst_mult_130_U8 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n8, B => 
                           dam_demodulator_inst_mult_130_n47, CI => 
                           dam_demodulator_inst_mult_130_n32, CO => 
                           dam_demodulator_inst_mult_130_n7, S => 
                           dam_demodulator_inst_prod_q_id_2);
   dam_demodulator_inst_mult_130_U7 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n7, B => 
                           dam_demodulator_inst_mult_130_n30, CI => 
                           dam_demodulator_inst_mult_130_n28, CO => 
                           dam_demodulator_inst_mult_130_n6, S => 
                           dam_demodulator_inst_prod_q_id_3);
   dam_demodulator_inst_mult_130_U6 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n22, B => 
                           dam_demodulator_inst_mult_130_n24, CI => 
                           dam_demodulator_inst_mult_130_n6, CO => 
                           dam_demodulator_inst_mult_130_n5, S => 
                           dam_demodulator_inst_prod_q_id_4);
   dam_demodulator_inst_mult_130_U5 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n16, B => 
                           dam_demodulator_inst_mult_130_n21, CI => 
                           dam_demodulator_inst_mult_130_n5, CO => 
                           dam_demodulator_inst_mult_130_n4, S => 
                           dam_demodulator_inst_prod_q_id_5);
   dam_demodulator_inst_mult_130_U4 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n12, B => 
                           dam_demodulator_inst_mult_130_n15, CI => 
                           dam_demodulator_inst_mult_130_n4, CO => 
                           dam_demodulator_inst_mult_130_n3, S => 
                           dam_demodulator_inst_prod_q_id_6);
   dam_demodulator_inst_mult_130_U3 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n11, B => 
                           dam_demodulator_inst_mult_130_n10, CI => 
                           dam_demodulator_inst_mult_130_n3, CO => 
                           dam_demodulator_inst_mult_130_n2, S => 
                           dam_demodulator_inst_prod_q_id_7);
   dam_demodulator_inst_mult_130_U2 : ADFULD1 port map( A => 
                           dam_demodulator_inst_mult_130_n9, B => 
                           dam_demodulator_inst_mult_130_n33, CI => 
                           dam_demodulator_inst_mult_130_n2, CO => 
                           dam_demodulator_inst_mult_130_n1, S => 
                           dam_demodulator_inst_prod_q_id_8);
   dam_demodulator_inst_sub_132_U12 : NOR2M1D1 port map( A1 => 
                           dam_demodulator_inst_prod_i_qd_0, A2 => 
                           dam_demodulator_inst_prod_q_id_0, Z => 
                           dam_demodulator_inst_sub_132_n10);
   dam_demodulator_inst_sub_132_U11 : AND2D1 port map( A1 => 
                           dam_demodulator_inst_sub_132_n10, A2 => 
                           dam_demodulator_inst_sub_132_n9, Z => 
                           dam_demodulator_inst_sub_132_n11);
   dam_demodulator_inst_sub_132_U10 : OAI22D1 port map( A1 => 
                           dam_demodulator_inst_sub_132_n10, A2 => 
                           dam_demodulator_inst_sub_132_n9, B1 => 
                           dam_demodulator_inst_prod_i_qd_1, B2 => 
                           dam_demodulator_inst_sub_132_n11, Z => 
                           dam_demodulator_inst_sub_132_carry_2_port);
   dam_demodulator_inst_sub_132_U9 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_i_qd_9, Z => 
                           dam_demodulator_inst_sub_132_n1);
   dam_demodulator_inst_sub_132_U8 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_i_qd_8, Z => 
                           dam_demodulator_inst_sub_132_n2);
   dam_demodulator_inst_sub_132_U7 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_1, Z => 
                           dam_demodulator_inst_sub_132_n9);
   dam_demodulator_inst_sub_132_U6 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_i_qd_7, Z => 
                           dam_demodulator_inst_sub_132_n3);
   dam_demodulator_inst_sub_132_U5 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_i_qd_4, Z => 
                           dam_demodulator_inst_sub_132_n6);
   dam_demodulator_inst_sub_132_U4 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_i_qd_2, Z => 
                           dam_demodulator_inst_sub_132_n8);
   dam_demodulator_inst_sub_132_U3 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_i_qd_6, Z => 
                           dam_demodulator_inst_sub_132_n4);
   dam_demodulator_inst_sub_132_U2 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_i_qd_5, Z => 
                           dam_demodulator_inst_sub_132_n5);
   dam_demodulator_inst_sub_132_U1 : INVD1 port map( A => 
                           dam_demodulator_inst_prod_i_qd_3, Z => 
                           dam_demodulator_inst_sub_132_n7);
   dam_demodulator_inst_sub_132_U2_2 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_2, B => 
                           dam_demodulator_inst_sub_132_n8, CI => 
                           dam_demodulator_inst_sub_132_carry_2_port, CO => 
                           dam_demodulator_inst_sub_132_carry_3_port, S => 
                           dam_demodulator_inst_result_2_port);
   dam_demodulator_inst_sub_132_U2_3 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_3, B => 
                           dam_demodulator_inst_sub_132_n7, CI => 
                           dam_demodulator_inst_sub_132_carry_3_port, CO => 
                           dam_demodulator_inst_sub_132_carry_4_port, S => 
                           dam_demodulator_inst_result_3_port);
   dam_demodulator_inst_sub_132_U2_4 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_4, B => 
                           dam_demodulator_inst_sub_132_n6, CI => 
                           dam_demodulator_inst_sub_132_carry_4_port, CO => 
                           dam_demodulator_inst_sub_132_carry_5_port, S => 
                           dam_demodulator_inst_result_4_port);
   dam_demodulator_inst_sub_132_U2_5 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_5, B => 
                           dam_demodulator_inst_sub_132_n5, CI => 
                           dam_demodulator_inst_sub_132_carry_5_port, CO => 
                           dam_demodulator_inst_sub_132_carry_6_port, S => 
                           dam_demodulator_inst_result_5_port);
   dam_demodulator_inst_sub_132_U2_6 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_6, B => 
                           dam_demodulator_inst_sub_132_n4, CI => 
                           dam_demodulator_inst_sub_132_carry_6_port, CO => 
                           dam_demodulator_inst_sub_132_carry_7_port, S => 
                           dam_demodulator_inst_result_6_port);
   dam_demodulator_inst_sub_132_U2_7 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_7, B => 
                           dam_demodulator_inst_sub_132_n3, CI => 
                           dam_demodulator_inst_sub_132_carry_7_port, CO => 
                           dam_demodulator_inst_sub_132_carry_8_port, S => 
                           dam_demodulator_inst_result_7_port);
   dam_demodulator_inst_sub_132_U2_8 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_8, B => 
                           dam_demodulator_inst_sub_132_n2, CI => 
                           dam_demodulator_inst_sub_132_carry_8_port, CO => 
                           dam_demodulator_inst_sub_132_carry_9_port, S => 
                           dam_demodulator_inst_result_8_port);
   dam_demodulator_inst_sub_132_U2_9 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_9, B => 
                           dam_demodulator_inst_sub_132_n1, CI => 
                           dam_demodulator_inst_sub_132_carry_9_port, CO => 
                           dam_demodulator_inst_sub_132_carry_10_port, S => 
                           dam_demodulator_inst_result_9_port);
   dam_demodulator_inst_sub_132_U2_10 : ADFULD1 port map( A => 
                           dam_demodulator_inst_prod_q_id_9, B => 
                           dam_demodulator_inst_sub_132_n1, CI => 
                           dam_demodulator_inst_sub_132_carry_10_port, CO => 
                           dam_demodulator_inst_sub_132_n_1004, S => 
                           dam_demodulator_inst_result_10_port);
   sl_slicer_inst_U14 : AOI21D1 port map( A1 => sl_slicer_inst_n8, A2 => 
                           sl_slicer_inst_n7, B => 
                           sl_slicer_inst_sum0_1_2_3_8_port, Z => 
                           sl_slicer_inst_N1);
   sl_slicer_inst_U13 : NOR4D1 port map( A1 => sl_slicer_inst_sum0_1_2_3_7_port
                           , A2 => sl_slicer_inst_sum0_1_2_3_6_port, A3 => 
                           sl_slicer_inst_sum0_1_2_3_5_port, A4 => 
                           sl_slicer_inst_sum0_1_2_3_4_port, Z => 
                           sl_slicer_inst_n7);
   sl_slicer_inst_U12 : NOR4D1 port map( A1 => sl_slicer_inst_sum0_1_2_3_3_port
                           , A2 => sl_slicer_inst_sum0_1_2_3_2_port, A3 => 
                           sl_slicer_inst_sum0_1_2_3_1_port, A4 => 
                           sl_slicer_inst_sum0_1_2_3_0_port, Z => 
                           sl_slicer_inst_n8);
   sl_slicer_inst_U11 : TIELO port map( Z => sl_slicer_inst_n101);
   sl_slicer_inst_U10 : INVD1 port map( A => clk4, Z => sl_slicer_inst_n6);
   sl_slicer_inst_U9 : INVD1 port map( A => 
                           sl_slicer_inst_arx_counter_reg_0_port, Z => 
                           sl_slicer_inst_n9);
   sl_slicer_inst_U3 : INVD1 port map( A => sl_slicer_inst_n6, Z => 
                           sl_slicer_inst_n100);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_1_6 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_20_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_13_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_0_6 : DFFRPQ1 port map( D => 
                           demodulator_out_6_port, CK => sl_slicer_inst_n100, 
                           RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_20_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_2_6 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_13_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_6_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_0_0 : DFFRPQ1 port map( D => 
                           demodulator_out_0_port, CK => sl_slicer_inst_n100, 
                           RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_14_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_1_1 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_15_port, CK => 
                           clk4, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_8_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_1_2 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_16_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_9_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_1_3 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_17_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_10_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_1_4 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_18_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_11_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_1_5 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_19_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_12_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_0_1 : DFFRPQ1 port map( D => 
                           demodulator_out_1_port, CK => sl_slicer_inst_n100, 
                           RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_15_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_0_2 : DFFRPQ1 port map( D => 
                           demodulator_out_2_port, CK => sl_slicer_inst_n100, 
                           RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_16_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_0_3 : DFFRPQ1 port map( D => 
                           demodulator_out_3_port, CK => sl_slicer_inst_n100, 
                           RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_17_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_0_4 : DFFRPQ1 port map( D => 
                           demodulator_out_4_port, CK => sl_slicer_inst_n100, 
                           RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_18_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_0_5 : DFFRPQ1 port map( D => 
                           demodulator_out_5_port, CK => sl_slicer_inst_n100, 
                           RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_19_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_1_0 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_14_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_7_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_2_0 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_7_port, CK => 
                           clk4, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_0_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_2_1 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_8_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_1_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_2_2 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_9_port, CK => 
                           clk4, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_2_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_2_3 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_10_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_3_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_2_4 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_11_port, CK => 
                           clk4, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_4_port);
   sl_slicer_inst_arx_slicer_fifo_reg_reg_2_5 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_arx_slicer_fifo_reg_12_port, CK => 
                           sl_slicer_inst_n100, RB => rstn, Q => 
                           sl_slicer_inst_arx_slicer_fifo_reg_5_port);
   sl_slicer_inst_arx_counter_reg_reg_1 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_counter_1, CK => clk4, RB => rstn, Q 
                           => sl_slicer_inst_arx_counter_reg_1_port);
   sl_slicer_inst_arx_counter_reg_reg_0 : DFFRPQ1 port map( D => 
                           sl_slicer_inst_n9, CK => sl_slicer_inst_n100, RB => 
                           rstn, Q => sl_slicer_inst_arx_counter_reg_0_port);
   sl_slicer_inst_arx_output_reg_reg : DFFRPQ1 port map( D => sl_slicer_inst_n5
                           , CK => clk4, RB => rstn, Q => slicer_out_port);
   sl_slicer_inst_U8 : EXNOR2D1 port map( A1 => 
                           sl_slicer_inst_arx_counter_reg_1_port, A2 => 
                           sl_slicer_inst_n9, Z => sl_slicer_inst_counter_1);
   sl_slicer_inst_U7 : EXOR2D1 port map( A1 => 
                           sl_slicer_inst_arx_counter_reg_1_port, A2 => 
                           n_Logic1, Z => sl_slicer_inst_n2);
   sl_slicer_inst_U6 : EXNOR2D1 port map( A1 => sl_slicer_inst_n9, A2 => 
                           n_Logic1, Z => sl_slicer_inst_n3);
   sl_slicer_inst_U5 : OAI21D1 port map( A1 => sl_slicer_inst_n2, A2 => 
                           sl_slicer_inst_n3, B => slicer_out_port, Z => 
                           sl_slicer_inst_n4);
   sl_slicer_inst_U4 : OAI31M10D1 port map( A1 => sl_slicer_inst_N1, A2 => 
                           sl_slicer_inst_n2, A3 => sl_slicer_inst_n3, B => 
                           sl_slicer_inst_n4, Z => sl_slicer_inst_n5);
   sl_slicer_inst_add_2_root_add_122_U2 : EXOR2D1 port map( A1 => 
                           sl_slicer_inst_arx_slicer_fifo_reg_14_port, A2 => 
                           demodulator_out_0_port, Z => sl_slicer_inst_sum2_3_0
                           );
   sl_slicer_inst_add_2_root_add_122_U1 : AND2D1 port map( A1 => 
                           sl_slicer_inst_arx_slicer_fifo_reg_14_port, A2 => 
                           demodulator_out_0_port, Z => 
                           sl_slicer_inst_add_2_root_add_122_n1);
   sl_slicer_inst_add_2_root_add_122_U1_1 : ADFULD1 port map( A => 
                           demodulator_out_1_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_15_port, CI => 
                           sl_slicer_inst_add_2_root_add_122_n1, CO => 
                           sl_slicer_inst_add_2_root_add_122_carry_2_port, S =>
                           sl_slicer_inst_sum2_3_1);
   sl_slicer_inst_add_2_root_add_122_U1_2 : ADFULD1 port map( A => 
                           demodulator_out_2_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_16_port, CI => 
                           sl_slicer_inst_add_2_root_add_122_carry_2_port, CO 
                           => sl_slicer_inst_add_2_root_add_122_carry_3_port, S
                           => sl_slicer_inst_sum2_3_2);
   sl_slicer_inst_add_2_root_add_122_U1_3 : ADFULD1 port map( A => 
                           demodulator_out_3_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_17_port, CI => 
                           sl_slicer_inst_add_2_root_add_122_carry_3_port, CO 
                           => sl_slicer_inst_add_2_root_add_122_carry_4_port, S
                           => sl_slicer_inst_sum2_3_3);
   sl_slicer_inst_add_2_root_add_122_U1_4 : ADFULD1 port map( A => 
                           demodulator_out_4_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_18_port, CI => 
                           sl_slicer_inst_add_2_root_add_122_carry_4_port, CO 
                           => sl_slicer_inst_add_2_root_add_122_carry_5_port, S
                           => sl_slicer_inst_sum2_3_4);
   sl_slicer_inst_add_2_root_add_122_U1_5 : ADFULD1 port map( A => 
                           demodulator_out_5_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_19_port, CI => 
                           sl_slicer_inst_add_2_root_add_122_carry_5_port, CO 
                           => sl_slicer_inst_add_2_root_add_122_carry_6_port, S
                           => sl_slicer_inst_sum2_3_5);
   sl_slicer_inst_add_2_root_add_122_U1_6 : ADFULD1 port map( A => 
                           demodulator_out_6_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_20_port, CI => 
                           sl_slicer_inst_add_2_root_add_122_carry_6_port, CO 
                           => sl_slicer_inst_add_2_root_add_122_carry_7_port, S
                           => sl_slicer_inst_sum2_3_6);
   sl_slicer_inst_add_2_root_add_122_U1_7 : ADFULD1 port map( A => 
                           demodulator_out_6_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_20_port, CI => 
                           sl_slicer_inst_add_2_root_add_122_carry_7_port, CO 
                           => sl_slicer_inst_add_2_root_add_122_n_1217, S => 
                           sl_slicer_inst_sum2_3_7);
   sl_slicer_inst_add_1_root_add_122_U2 : EXOR2D1 port map( A1 => 
                           sl_slicer_inst_arx_slicer_fifo_reg_0_port, A2 => 
                           sl_slicer_inst_arx_slicer_fifo_reg_7_port, Z => 
                           sl_slicer_inst_sum0_1_0);
   sl_slicer_inst_add_1_root_add_122_U1 : AND2D1 port map( A1 => 
                           sl_slicer_inst_arx_slicer_fifo_reg_0_port, A2 => 
                           sl_slicer_inst_arx_slicer_fifo_reg_7_port, Z => 
                           sl_slicer_inst_add_1_root_add_122_n1);
   sl_slicer_inst_add_1_root_add_122_U1_1 : ADFULD1 port map( A => 
                           sl_slicer_inst_arx_slicer_fifo_reg_8_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_1_port, CI => 
                           sl_slicer_inst_add_1_root_add_122_n1, CO => 
                           sl_slicer_inst_add_1_root_add_122_carry_2_port, S =>
                           sl_slicer_inst_sum0_1_1);
   sl_slicer_inst_add_1_root_add_122_U1_2 : ADFULD1 port map( A => 
                           sl_slicer_inst_arx_slicer_fifo_reg_9_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_2_port, CI => 
                           sl_slicer_inst_add_1_root_add_122_carry_2_port, CO 
                           => sl_slicer_inst_add_1_root_add_122_carry_3_port, S
                           => sl_slicer_inst_sum0_1_2);
   sl_slicer_inst_add_1_root_add_122_U1_3 : ADFULD1 port map( A => 
                           sl_slicer_inst_arx_slicer_fifo_reg_10_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_3_port, CI => 
                           sl_slicer_inst_add_1_root_add_122_carry_3_port, CO 
                           => sl_slicer_inst_add_1_root_add_122_carry_4_port, S
                           => sl_slicer_inst_sum0_1_3);
   sl_slicer_inst_add_1_root_add_122_U1_4 : ADFULD1 port map( A => 
                           sl_slicer_inst_arx_slicer_fifo_reg_11_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_4_port, CI => 
                           sl_slicer_inst_add_1_root_add_122_carry_4_port, CO 
                           => sl_slicer_inst_add_1_root_add_122_carry_5_port, S
                           => sl_slicer_inst_sum0_1_4);
   sl_slicer_inst_add_1_root_add_122_U1_5 : ADFULD1 port map( A => 
                           sl_slicer_inst_arx_slicer_fifo_reg_12_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_5_port, CI => 
                           sl_slicer_inst_add_1_root_add_122_carry_5_port, CO 
                           => sl_slicer_inst_add_1_root_add_122_carry_6_port, S
                           => sl_slicer_inst_sum0_1_5);
   sl_slicer_inst_add_1_root_add_122_U1_6 : ADFULD1 port map( A => 
                           sl_slicer_inst_arx_slicer_fifo_reg_13_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_6_port, CI => 
                           sl_slicer_inst_add_1_root_add_122_carry_6_port, CO 
                           => sl_slicer_inst_add_1_root_add_122_carry_7_port, S
                           => sl_slicer_inst_sum0_1_6);
   sl_slicer_inst_add_1_root_add_122_U1_7 : ADFULD1 port map( A => 
                           sl_slicer_inst_arx_slicer_fifo_reg_13_port, B => 
                           sl_slicer_inst_arx_slicer_fifo_reg_6_port, CI => 
                           sl_slicer_inst_add_1_root_add_122_carry_7_port, CO 
                           => sl_slicer_inst_add_1_root_add_122_n_1220, S => 
                           sl_slicer_inst_sum0_1_7);
   sl_slicer_inst_add_0_root_add_122_U2 : EXOR2D1 port map( A1 => 
                           sl_slicer_inst_sum0_1_0, A2 => 
                           sl_slicer_inst_sum2_3_0, Z => 
                           sl_slicer_inst_sum0_1_2_3_0_port);
   sl_slicer_inst_add_0_root_add_122_U1 : AND2D1 port map( A1 => 
                           sl_slicer_inst_sum0_1_0, A2 => 
                           sl_slicer_inst_sum2_3_0, Z => 
                           sl_slicer_inst_add_0_root_add_122_n1);
   sl_slicer_inst_add_0_root_add_122_U1_1 : ADFULD1 port map( A => 
                           sl_slicer_inst_sum2_3_1, B => 
                           sl_slicer_inst_sum0_1_1, CI => 
                           sl_slicer_inst_add_0_root_add_122_n1, CO => 
                           sl_slicer_inst_add_0_root_add_122_carry_2_port, S =>
                           sl_slicer_inst_sum0_1_2_3_1_port);
   sl_slicer_inst_add_0_root_add_122_U1_2 : ADFULD1 port map( A => 
                           sl_slicer_inst_sum2_3_2, B => 
                           sl_slicer_inst_sum0_1_2, CI => 
                           sl_slicer_inst_add_0_root_add_122_carry_2_port, CO 
                           => sl_slicer_inst_add_0_root_add_122_carry_3_port, S
                           => sl_slicer_inst_sum0_1_2_3_2_port);
   sl_slicer_inst_add_0_root_add_122_U1_3 : ADFULD1 port map( A => 
                           sl_slicer_inst_sum2_3_3, B => 
                           sl_slicer_inst_sum0_1_3, CI => 
                           sl_slicer_inst_add_0_root_add_122_carry_3_port, CO 
                           => sl_slicer_inst_add_0_root_add_122_carry_4_port, S
                           => sl_slicer_inst_sum0_1_2_3_3_port);
   sl_slicer_inst_add_0_root_add_122_U1_4 : ADFULD1 port map( A => 
                           sl_slicer_inst_sum2_3_4, B => 
                           sl_slicer_inst_sum0_1_4, CI => 
                           sl_slicer_inst_add_0_root_add_122_carry_4_port, CO 
                           => sl_slicer_inst_add_0_root_add_122_carry_5_port, S
                           => sl_slicer_inst_sum0_1_2_3_4_port);
   sl_slicer_inst_add_0_root_add_122_U1_5 : ADFULD1 port map( A => 
                           sl_slicer_inst_sum2_3_5, B => 
                           sl_slicer_inst_sum0_1_5, CI => 
                           sl_slicer_inst_add_0_root_add_122_carry_5_port, CO 
                           => sl_slicer_inst_add_0_root_add_122_carry_6_port, S
                           => sl_slicer_inst_sum0_1_2_3_5_port);
   sl_slicer_inst_add_0_root_add_122_U1_6 : ADFULD1 port map( A => 
                           sl_slicer_inst_sum2_3_6, B => 
                           sl_slicer_inst_sum0_1_6, CI => 
                           sl_slicer_inst_add_0_root_add_122_carry_6_port, CO 
                           => sl_slicer_inst_add_0_root_add_122_carry_7_port, S
                           => sl_slicer_inst_sum0_1_2_3_6_port);
   sl_slicer_inst_add_0_root_add_122_U1_7 : ADFULD1 port map( A => 
                           sl_slicer_inst_sum2_3_7, B => 
                           sl_slicer_inst_sum0_1_7, CI => 
                           sl_slicer_inst_add_0_root_add_122_carry_7_port, CO 
                           => sl_slicer_inst_add_0_root_add_122_carry_8_port, S
                           => sl_slicer_inst_sum0_1_2_3_7_port);
   sl_slicer_inst_add_0_root_add_122_U1_8 : ADFULD1 port map( A => 
                           sl_slicer_inst_sum2_3_7, B => 
                           sl_slicer_inst_sum0_1_7, CI => 
                           sl_slicer_inst_add_0_root_add_122_carry_8_port, CO 
                           => sl_slicer_inst_add_0_root_add_122_n_1223, S => 
                           sl_slicer_inst_sum0_1_2_3_8_port);

end flat_structure_none_10;
