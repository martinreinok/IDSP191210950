
library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

package CONV_PACK_sec_df2_std is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_sec_df2_std;

library IEEE,umcl18u250t2;

use IEEE.std_logic_1164.all;
use umcl18u250t2.umcl18u250t2_VCOMPONENTS.all;

use work.CONV_PACK_sec_df2_std.all;

architecture flat_rtl_none_10 of sec_df2_std is

   component ADFULD1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component EXOR3D1
      port( A1, A2, A3 : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21M20D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21D1
      port( A1, A2, B : in std_logic;  Z : out std_logic);
   end component;
   
   component ADHALFDL
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component INVD1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component EXOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  Z : out std_logic);
   end component;
   
   component NAN2M1D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFRPQ1
      port( D, CK, RB : in std_logic;  Q : out std_logic);
   end component;
   
   component TIEHI
      port( Z : out std_logic);
   end component;
   
   component TIELO
      port( Z : out std_logic);
   end component;
   
   signal sec_df2_inst_n_1064, sec_df2_inst_n_1063, sec_df2_inst_n_1062, 
      sec_df2_inst_n_1061, sec_df2_inst_n_1060, sec_df2_inst_n_1059, 
      sec_df2_inst_n_1058, sec_df2_inst_n_1057, sec_df2_inst_n_1056, 
      sec_df2_inst_n_1055, sec_df2_inst_n_1054, sec_df2_inst_n_1053, 
      sec_df2_inst_n_1052, sec_df2_inst_n_1051, sec_df2_inst_n_1050, 
      sec_df2_inst_n_1049, sec_df2_inst_n_1048, sec_df2_inst_n_1047, 
      sec_df2_inst_n_1046, sec_df2_inst_n_1045, sec_df2_inst_n_1044, 
      sec_df2_inst_n_1043, sec_df2_inst_n_1042, sec_df2_inst_n_1041, 
      sec_df2_inst_n90, sec_df2_inst_n80, sec_df2_inst_n70, sec_df2_inst_n60, 
      sec_df2_inst_n50, sec_df2_inst_n40, sec_df2_inst_n30, sec_df2_inst_n27, 
      sec_df2_inst_n110, sec_df2_inst_add_416_C138_rn_carry_7_port, 
      sec_df2_inst_add_416_C138_rn_carry_6_port, 
      sec_df2_inst_add_416_C138_rn_carry_5_port, 
      sec_df2_inst_add_416_C138_rn_carry_4_port, 
      sec_df2_inst_add_416_C138_rn_carry_3_port, 
      sec_df2_inst_add_416_C138_rn_carry_2_port, 
      sec_df2_inst_add_416_C138_rn_carry_1_port, 
      sec_df2_inst_add_139_carry_14_port, sec_df2_inst_add_139_carry_13_port, 
      sec_df2_inst_add_139_carry_12_port, sec_df2_inst_add_139_carry_11_port, 
      sec_df2_inst_add_139_carry_10_port, sec_df2_inst_add_139_carry_9_port, 
      sec_df2_inst_add_139_carry_8_port, sec_df2_inst_mult_133_n1, 
      sec_df2_inst_mult_133_n2, sec_df2_inst_mult_133_n3, 
      sec_df2_inst_mult_133_n4, sec_df2_inst_mult_133_n5, 
      sec_df2_inst_mult_133_n6, sec_df2_inst_mult_133_n7, 
      sec_df2_inst_mult_133_n8, sec_df2_inst_mult_133_n9, 
      sec_df2_inst_mult_133_n10, sec_df2_inst_mult_133_n11, 
      sec_df2_inst_mult_133_n12, sec_df2_inst_mult_133_n13, 
      sec_df2_inst_mult_133_n15, sec_df2_inst_mult_133_n16, 
      sec_df2_inst_mult_133_n17, sec_df2_inst_mult_133_n18, 
      sec_df2_inst_mult_133_n19, sec_df2_inst_mult_133_n20, 
      sec_df2_inst_mult_133_n21, sec_df2_inst_mult_133_n22, 
      sec_df2_inst_mult_133_n23, sec_df2_inst_mult_133_n24, 
      sec_df2_inst_mult_133_n25, sec_df2_inst_mult_133_n26, 
      sec_df2_inst_mult_131_n2, sec_df2_inst_mult_131_n3, 
      sec_df2_inst_mult_131_n4, sec_df2_inst_mult_131_n5, 
      sec_df2_inst_mult_131_n6, sec_df2_inst_mult_131_n7, 
      sec_df2_inst_mult_131_n8, sec_df2_inst_mult_131_n9, 
      sec_df2_inst_mult_131_n10, sec_df2_inst_mult_131_n11, 
      sec_df2_inst_mult_131_n12, sec_df2_inst_mult_131_n13, 
      sec_df2_inst_mult_131_n14, sec_df2_inst_mult_131_n15, 
      sec_df2_inst_mult_131_n16, sec_df2_inst_mult_134_n1, 
      sec_df2_inst_mult_134_n2, sec_df2_inst_mult_134_n3, 
      sec_df2_inst_mult_134_n4, sec_df2_inst_mult_134_n5, 
      sec_df2_inst_mult_134_n6, sec_df2_inst_mult_134_n7, 
      sec_df2_inst_mult_134_n8, sec_df2_inst_mult_134_n9, 
      sec_df2_inst_mult_134_n10, sec_df2_inst_mult_134_n11, 
      sec_df2_inst_mult_134_n16, sec_df2_inst_mult_134_n17, 
      sec_df2_inst_mult_134_n18, sec_df2_inst_mult_134_n19, 
      sec_df2_inst_mult_134_n20, sec_df2_inst_mult_134_n21, 
      sec_df2_inst_mult_134_n22, sec_df2_inst_mult_134_n23, 
      sec_df2_inst_mult_134_n24, sec_df2_inst_mult_134_n25, 
      sec_df2_inst_add_416_C139_rn_carry_7_port, 
      sec_df2_inst_add_416_C139_rn_carry_6_port, 
      sec_df2_inst_add_416_C139_rn_carry_5_port, 
      sec_df2_inst_add_416_C139_rn_carry_4_port, 
      sec_df2_inst_add_416_C139_rn_carry_3_port, 
      sec_df2_inst_add_416_C139_rn_carry_2_port, 
      sec_df2_inst_add_416_C139_rn_carry_1_port, sec_df2_inst_m3_0, 
      sec_df2_inst_m3_10, sec_df2_inst_m3_11, sec_df2_inst_m3_12, 
      sec_df2_inst_m3_13, sec_df2_inst_m3_14, sec_df2_inst_m3_1, 
      sec_df2_inst_m3_2, sec_df2_inst_m3_3, sec_df2_inst_m3_4, 
      sec_df2_inst_m3_5, sec_df2_inst_m3_6, sec_df2_inst_m3_7, 
      sec_df2_inst_m3_8, sec_df2_inst_m3_9, sec_df2_inst_m5_10, 
      sec_df2_inst_m5_11, sec_df2_inst_m5_12, sec_df2_inst_m5_13, 
      sec_df2_inst_m5_1, sec_df2_inst_m5_2, sec_df2_inst_m5_3, 
      sec_df2_inst_m5_4, sec_df2_inst_m5_5, sec_df2_inst_m5_6, 
      sec_df2_inst_m5_7, sec_df2_inst_m5_8, sec_df2_inst_m5_9, 
      sec_df2_inst_m5_15, sec_df2_inst_m2_10, sec_df2_inst_m2_11, 
      sec_df2_inst_m2_12, sec_df2_inst_m2_13, sec_df2_inst_m2_14, 
      sec_df2_inst_m2_1, sec_df2_inst_m2_2, sec_df2_inst_m2_3, 
      sec_df2_inst_m2_4, sec_df2_inst_m2_5, sec_df2_inst_m2_6, 
      sec_df2_inst_m2_7, sec_df2_inst_m2_8, sec_df2_inst_m2_9, 
      sec_df2_inst_m4_0, sec_df2_inst_m4_10, sec_df2_inst_m4_11, 
      sec_df2_inst_m4_12, sec_df2_inst_m4_13, sec_df2_inst_m4_1, 
      sec_df2_inst_m4_2, sec_df2_inst_m4_3, sec_df2_inst_m4_4, 
      sec_df2_inst_m4_5, sec_df2_inst_m4_6, sec_df2_inst_m4_7, 
      sec_df2_inst_m4_8, sec_df2_inst_m4_9, sec_df2_inst_m4_15, 
      sec_df2_inst_m1_10, sec_df2_inst_m1_11, sec_df2_inst_m1_12, 
      sec_df2_inst_m1_13, sec_df2_inst_m1_7, sec_df2_inst_m1_8, 
      sec_df2_inst_m1_9, sec_df2_inst_m1_15, sec_df2_inst_p4_0, 
      sec_df2_inst_p4_1, sec_df2_inst_p4_2, sec_df2_inst_p4_3, 
      sec_df2_inst_p4_4, sec_df2_inst_p4_5, sec_df2_inst_p4_6, 
      sec_df2_inst_p4_7, sec_df2_inst_N26, sec_df2_inst_N25, sec_df2_inst_N24, 
      sec_df2_inst_N23, sec_df2_inst_N22, sec_df2_inst_N21, sec_df2_inst_N20, 
      sec_df2_inst_N19, sec_df2_inst_N18, sec_df2_inst_N17, sec_df2_inst_N16, 
      sec_df2_inst_N15, sec_df2_inst_N14, sec_df2_inst_N13, sec_df2_inst_N12, 
      sec_df2_inst_N11, sec_df2_inst_N10, sec_df2_inst_N9, sec_df2_inst_N8, 
      sec_df2_inst_N7, sec_df2_inst_N6, sec_df2_inst_N5, sec_df2_inst_N4, 
      sec_df2_inst_N3, sec_df2_inst_N2, sec_df2_inst_N1, sec_df2_inst_N0, 
      sec_df2_inst_p2_0_port, sec_df2_inst_p2_1_port, sec_df2_inst_p2_2_port, 
      sec_df2_inst_p2_3_port, sec_df2_inst_p2_4_port, sec_df2_inst_p2_5_port, 
      sec_df2_inst_p2_6_port, sec_df2_inst_p2_7_port, sec_df2_inst_p1_0_port, 
      sec_df2_inst_p1_1_port, sec_df2_inst_p1_2_port, sec_df2_inst_p1_3_port, 
      sec_df2_inst_p1_4_port, sec_df2_inst_p1_5_port, sec_df2_inst_p1_6_port, 
      sec_df2_inst_p1_7_port, sec_df2_inst_arx_z2_reg_3_port, 
      sec_df2_inst_arx_z2_reg_4_port, sec_df2_inst_arx_z2_reg_5_port, 
      sec_df2_inst_arx_z2_reg_6_port, sec_df2_inst_arx_z2_reg_7_port, 
      sec_df2_inst_arx_z1_reg_2_port, sec_df2_inst_arx_z1_reg_3_port, 
      sec_df2_inst_arx_z1_reg_4_port, sec_df2_inst_arx_z1_reg_5_port, 
      sec_df2_inst_arx_z1_reg_6_port, 
      sec_df2_inst_add_1_root_add_136_carry_1_port, 
      sec_df2_inst_add_1_root_add_136_carry_2_port, 
      sec_df2_inst_add_1_root_add_136_carry_3_port, 
      sec_df2_inst_add_1_root_add_136_carry_4_port, 
      sec_df2_inst_add_1_root_add_136_carry_5_port, 
      sec_df2_inst_add_1_root_add_136_carry_6_port, 
      sec_df2_inst_add_1_root_add_136_carry_7_port, sec_df2_inst_mult_137_n78, 
      sec_df2_inst_mult_137_n77, sec_df2_inst_mult_137_n76, 
      sec_df2_inst_mult_137_n75, sec_df2_inst_mult_137_n74, 
      sec_df2_inst_mult_137_n73, sec_df2_inst_mult_137_n72, 
      sec_df2_inst_mult_137_n71, sec_df2_inst_mult_137_n70, 
      sec_df2_inst_mult_137_n69, sec_df2_inst_mult_137_n68, 
      sec_df2_inst_mult_137_n25, sec_df2_inst_mult_137_n24, 
      sec_df2_inst_mult_137_n23, sec_df2_inst_mult_137_n22, 
      sec_df2_inst_mult_137_n21, sec_df2_inst_mult_137_n20, 
      sec_df2_inst_mult_137_n19, sec_df2_inst_mult_137_n18, 
      sec_df2_inst_mult_137_n17, sec_df2_inst_mult_137_n16, 
      sec_df2_inst_mult_137_n9, sec_df2_inst_mult_137_n8, 
      sec_df2_inst_mult_137_n7, sec_df2_inst_mult_137_n6, 
      sec_df2_inst_mult_137_n5, sec_df2_inst_mult_137_n4, 
      sec_df2_inst_mult_137_n3, sec_df2_inst_mult_137_n2, 
      sec_df2_inst_mult_137_n1, sec_df2_inst_add_135_n9, 
      sec_df2_inst_add_135_n8, sec_df2_inst_add_135_n7, sec_df2_inst_add_135_n6
      , sec_df2_inst_add_135_n5, sec_df2_inst_add_135_n4, 
      sec_df2_inst_add_135_n3, sec_df2_inst_add_135_n2, sec_df2_inst_add_135_n1
      , sec_df2_inst_add_135_carry_6_port, sec_df2_inst_add_135_carry_7_port, 
      sec_df2_inst_add_135_carry_8_port, sec_df2_inst_add_135_carry_9_port, 
      sec_df2_inst_add_135_carry_10_port, sec_df2_inst_add_135_carry_11_port, 
      sec_df2_inst_add_135_carry_12_port, sec_df2_inst_add_135_carry_13_port, 
      sec_df2_inst_add_135_carry_14_port, sec_df2_inst_mult_132_n89, 
      sec_df2_inst_mult_132_n88, sec_df2_inst_mult_132_n87, 
      sec_df2_inst_mult_132_n86, sec_df2_inst_mult_132_n85, 
      sec_df2_inst_mult_132_n84, sec_df2_inst_mult_132_n83, 
      sec_df2_inst_mult_132_n36, sec_df2_inst_mult_132_n35, 
      sec_df2_inst_mult_132_n34, sec_df2_inst_mult_132_n33, 
      sec_df2_inst_mult_132_n32, sec_df2_inst_mult_132_n31, 
      sec_df2_inst_mult_132_n30, sec_df2_inst_mult_132_n29, 
      sec_df2_inst_mult_132_n28, sec_df2_inst_mult_132_n27, 
      sec_df2_inst_mult_132_n26, sec_df2_inst_mult_132_n25, 
      sec_df2_inst_mult_132_n24, sec_df2_inst_mult_132_n23, 
      sec_df2_inst_mult_132_n22, sec_df2_inst_mult_132_n21, 
      sec_df2_inst_mult_132_n20, sec_df2_inst_mult_132_n19, 
      sec_df2_inst_mult_132_n18, sec_df2_inst_mult_132_n17, 
      sec_df2_inst_mult_132_n16, sec_df2_inst_mult_132_n15, 
      sec_df2_inst_mult_132_n14, sec_df2_inst_mult_132_n13, 
      sec_df2_inst_mult_132_n12, sec_df2_inst_mult_132_n11, 
      sec_df2_inst_mult_132_n10, sec_df2_inst_mult_132_n9, 
      sec_df2_inst_mult_132_n8, sec_df2_inst_mult_132_n7, 
      sec_df2_inst_mult_132_n6, sec_df2_inst_mult_132_n5, 
      sec_df2_inst_mult_132_n4, sec_df2_inst_mult_132_n3, 
      sec_df2_inst_mult_132_n2, sec_df2_inst_add_138_n8, 
      sec_df2_inst_add_138_n7, sec_df2_inst_add_138_n6, sec_df2_inst_add_138_n5
      , sec_df2_inst_add_138_n4, sec_df2_inst_add_138_n3, 
      sec_df2_inst_add_138_n2, sec_df2_inst_add_138_n1, 
      sec_df2_inst_add_138_carry_6_port, sec_df2_inst_add_138_carry_7_port, 
      sec_df2_inst_add_138_carry_8_port, sec_df2_inst_add_138_carry_9_port, 
      sec_df2_inst_add_138_carry_10_port, sec_df2_inst_add_138_carry_11_port, 
      sec_df2_inst_add_138_carry_12_port, sec_df2_inst_add_138_carry_13_port, 
      sec_df2_inst_add_138_carry_14_port : std_logic;

begin
   
   sec_df2_inst_U50 : EXOR2D1 port map( A1 => sec_df2_inst_arx_z2_reg_3_port, 
                           A2 => sec_df2_inst_m4_0, Z => sec_df2_inst_m5_3);
   sec_df2_inst_U49 : NAN2D1 port map( A1 => sec_df2_inst_m4_0, A2 => 
                           sec_df2_inst_n40, Z => sec_df2_inst_mult_134_n11);
   sec_df2_inst_U48 : EXOR2D1 port map( A1 => sec_df2_inst_n70, A2 => 
                           sec_df2_inst_m4_0, Z => sec_df2_inst_mult_133_n26);
   sec_df2_inst_U47 : NAN2D1 port map( A1 => sec_df2_inst_m4_0, A2 => 
                           sec_df2_inst_arx_z2_reg_6_port, Z => 
                           sec_df2_inst_mult_133_n25);
   sec_df2_inst_U46 : EXOR2D1 port map( A1 => sec_df2_inst_N9, A2 => 
                           sec_df2_inst_N10, Z => sec_df2_inst_p4_0);
   sec_df2_inst_U45 : AND2D1 port map( A1 => sec_df2_inst_N9, A2 => 
                           sec_df2_inst_N10, Z => 
                           sec_df2_inst_add_416_C138_rn_carry_1_port);
   sec_df2_inst_U44 : EXOR2D1 port map( A1 => sec_df2_inst_N11, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_1_port, Z => 
                           sec_df2_inst_p4_1);
   sec_df2_inst_U43 : AND2D1 port map( A1 => sec_df2_inst_N11, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_1_port, Z => 
                           sec_df2_inst_add_416_C138_rn_carry_2_port);
   sec_df2_inst_U42 : EXOR2D1 port map( A1 => sec_df2_inst_N12, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_2_port, Z => 
                           sec_df2_inst_p4_2);
   sec_df2_inst_U41 : AND2D1 port map( A1 => sec_df2_inst_N12, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_2_port, Z => 
                           sec_df2_inst_add_416_C138_rn_carry_3_port);
   sec_df2_inst_U40 : EXOR2D1 port map( A1 => sec_df2_inst_N13, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_3_port, Z => 
                           sec_df2_inst_p4_3);
   sec_df2_inst_U39 : AND2D1 port map( A1 => sec_df2_inst_N13, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_3_port, Z => 
                           sec_df2_inst_add_416_C138_rn_carry_4_port);
   sec_df2_inst_U38 : EXOR2D1 port map( A1 => sec_df2_inst_N14, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_4_port, Z => 
                           sec_df2_inst_p4_4);
   sec_df2_inst_U37 : AND2D1 port map( A1 => sec_df2_inst_N14, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_4_port, Z => 
                           sec_df2_inst_add_416_C138_rn_carry_5_port);
   sec_df2_inst_U36 : EXOR2D1 port map( A1 => sec_df2_inst_N15, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_5_port, Z => 
                           sec_df2_inst_p4_5);
   sec_df2_inst_U35 : AND2D1 port map( A1 => sec_df2_inst_N15, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_5_port, Z => 
                           sec_df2_inst_add_416_C138_rn_carry_6_port);
   sec_df2_inst_U34 : EXOR2D1 port map( A1 => sec_df2_inst_N16, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_6_port, Z => 
                           sec_df2_inst_p4_6);
   sec_df2_inst_U33 : AND2D1 port map( A1 => sec_df2_inst_N16, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_6_port, Z => 
                           sec_df2_inst_add_416_C138_rn_carry_7_port);
   sec_df2_inst_U32 : EXOR2D1 port map( A1 => sec_df2_inst_N17, A2 => 
                           sec_df2_inst_add_416_C138_rn_carry_7_port, Z => 
                           sec_df2_inst_p4_7);
   sec_df2_inst_U31 : EXOR2D1 port map( A1 => sec_df2_inst_p4_0, A2 => 
                           sec_df2_inst_m1_7, Z => sec_df2_inst_N19);
   sec_df2_inst_U30 : AND2D1 port map( A1 => sec_df2_inst_m1_7, A2 => 
                           sec_df2_inst_p4_0, Z => 
                           sec_df2_inst_add_139_carry_8_port);
   sec_df2_inst_U29 : EXOR2D1 port map( A1 => sec_df2_inst_N18, A2 => 
                           sec_df2_inst_N19, Z => sec_df2_inst_p2_0_port);
   sec_df2_inst_U28 : AND2D1 port map( A1 => sec_df2_inst_N18, A2 => 
                           sec_df2_inst_N19, Z => 
                           sec_df2_inst_add_416_C139_rn_carry_1_port);
   sec_df2_inst_U27 : EXOR2D1 port map( A1 => sec_df2_inst_N20, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_1_port, Z => 
                           sec_df2_inst_p2_1_port);
   sec_df2_inst_U26 : AND2D1 port map( A1 => sec_df2_inst_N20, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_1_port, Z => 
                           sec_df2_inst_add_416_C139_rn_carry_2_port);
   sec_df2_inst_U25 : EXOR2D1 port map( A1 => sec_df2_inst_N21, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_2_port, Z => 
                           sec_df2_inst_p2_2_port);
   sec_df2_inst_U24 : AND2D1 port map( A1 => sec_df2_inst_N21, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_2_port, Z => 
                           sec_df2_inst_add_416_C139_rn_carry_3_port);
   sec_df2_inst_U23 : EXOR2D1 port map( A1 => sec_df2_inst_N22, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_3_port, Z => 
                           sec_df2_inst_p2_3_port);
   sec_df2_inst_U22 : AND2D1 port map( A1 => sec_df2_inst_N22, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_3_port, Z => 
                           sec_df2_inst_add_416_C139_rn_carry_4_port);
   sec_df2_inst_U21 : EXOR2D1 port map( A1 => sec_df2_inst_N23, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_4_port, Z => 
                           sec_df2_inst_p2_4_port);
   sec_df2_inst_U20 : AND2D1 port map( A1 => sec_df2_inst_N23, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_4_port, Z => 
                           sec_df2_inst_add_416_C139_rn_carry_5_port);
   sec_df2_inst_U19 : EXOR2D1 port map( A1 => sec_df2_inst_N24, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_5_port, Z => 
                           sec_df2_inst_p2_5_port);
   sec_df2_inst_U18 : AND2D1 port map( A1 => sec_df2_inst_N24, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_5_port, Z => 
                           sec_df2_inst_add_416_C139_rn_carry_6_port);
   sec_df2_inst_U17 : EXOR2D1 port map( A1 => sec_df2_inst_N25, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_6_port, Z => 
                           sec_df2_inst_p2_6_port);
   sec_df2_inst_U16 : AND2D1 port map( A1 => sec_df2_inst_N25, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_6_port, Z => 
                           sec_df2_inst_add_416_C139_rn_carry_7_port);
   sec_df2_inst_U15 : EXOR2D1 port map( A1 => sec_df2_inst_N26, A2 => 
                           sec_df2_inst_add_416_C139_rn_carry_7_port, Z => 
                           sec_df2_inst_p2_7_port);
   sec_df2_inst_U14 : TIELO port map( Z => sec_df2_inst_m3_0);
   sec_df2_inst_U13 : TIEHI port map( Z => sec_df2_inst_n90);
   sec_df2_inst_U12 : INVD1 port map( A => sec_df2_inst_mult_134_n1, Z => 
                           sec_df2_inst_m5_15);
   sec_df2_inst_U11 : INVD1 port map( A => sec_df2_inst_arx_z2_reg_7_port, Z =>
                           sec_df2_inst_n80);
   sec_df2_inst_U10 : INVD1 port map( A => sec_df2_inst_arx_z2_reg_5_port, Z =>
                           sec_df2_inst_n60);
   sec_df2_inst_U9 : INVD1 port map( A => sec_df2_inst_arx_z2_reg_6_port, Z => 
                           sec_df2_inst_n70);
   sec_df2_inst_U8 : INVD1 port map( A => sec_df2_inst_arx_z2_reg_4_port, Z => 
                           sec_df2_inst_n50);
   sec_df2_inst_U7 : INVD1 port map( A => sec_df2_inst_arx_z2_reg_3_port, Z => 
                           sec_df2_inst_n40);
   sec_df2_inst_U6 : INVD1 port map( A => sec_df2_inst_m5_2, Z => 
                           sec_df2_inst_n30);
   sec_df2_inst_U5 : INVD1 port map( A => sec_df2_inst_m5_1, Z => 
                           sec_df2_inst_n27);
   sec_df2_inst_U4 : INVD1 port map( A => sec_df2_inst_m4_0, Z => 
                           sec_df2_inst_n110);
   sec_df2_inst_U3 : INVD1 port map( A => sec_df2_inst_mult_133_n1, Z => 
                           sec_df2_inst_m4_15);
   sec_df2_inst_arx_p2_out_reg_reg_0 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p2_0_port, CK => clock, RB => resetn, Q
                           => data_out(0));
   sec_df2_inst_arx_p2_out_reg_reg_1 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p2_1_port, CK => clock, RB => resetn, Q
                           => data_out(1));
   sec_df2_inst_arx_p2_out_reg_reg_2 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p2_2_port, CK => clock, RB => resetn, Q
                           => data_out(2));
   sec_df2_inst_arx_p2_out_reg_reg_3 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p2_3_port, CK => clock, RB => resetn, Q
                           => data_out(3));
   sec_df2_inst_arx_p2_out_reg_reg_4 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p2_4_port, CK => clock, RB => resetn, Q
                           => data_out(4));
   sec_df2_inst_arx_p2_out_reg_reg_5 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p2_5_port, CK => clock, RB => resetn, Q
                           => data_out(5));
   sec_df2_inst_arx_p2_out_reg_reg_6 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p2_6_port, CK => clock, RB => resetn, Q
                           => data_out(6));
   sec_df2_inst_arx_p2_out_reg_reg_7 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p2_7_port, CK => clock, RB => resetn, Q
                           => data_out(7));
   sec_df2_inst_arx_z1_reg_reg_1 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p1_1_port, CK => clock, RB => resetn, Q
                           => sec_df2_inst_m3_2);
   sec_df2_inst_arx_z1_reg_reg_0 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p1_0_port, CK => clock, RB => resetn, Q
                           => sec_df2_inst_m3_1);
   sec_df2_inst_arx_z2_reg_reg_1 : DFFRPQ1 port map( D => sec_df2_inst_m3_2, CK
                           => clock, RB => resetn, Q => sec_df2_inst_m5_1);
   sec_df2_inst_arx_z2_reg_reg_0 : DFFRPQ1 port map( D => sec_df2_inst_m3_1, CK
                           => clock, RB => resetn, Q => sec_df2_inst_m4_0);
   sec_df2_inst_arx_z1_reg_reg_2 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p1_2_port, CK => clock, RB => resetn, Q
                           => sec_df2_inst_arx_z1_reg_2_port);
   sec_df2_inst_arx_z2_reg_reg_2 : DFFRPQ1 port map( D => 
                           sec_df2_inst_arx_z1_reg_2_port, CK => clock, RB => 
                           resetn, Q => sec_df2_inst_m5_2);
   sec_df2_inst_arx_z1_reg_reg_3 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p1_3_port, CK => clock, RB => resetn, Q
                           => sec_df2_inst_arx_z1_reg_3_port);
   sec_df2_inst_arx_z2_reg_reg_3 : DFFRPQ1 port map( D => 
                           sec_df2_inst_arx_z1_reg_3_port, CK => clock, RB => 
                           resetn, Q => sec_df2_inst_arx_z2_reg_3_port);
   sec_df2_inst_arx_z2_reg_reg_4 : DFFRPQ1 port map( D => 
                           sec_df2_inst_arx_z1_reg_4_port, CK => clock, RB => 
                           resetn, Q => sec_df2_inst_arx_z2_reg_4_port);
   sec_df2_inst_arx_z1_reg_reg_4 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p1_4_port, CK => clock, RB => resetn, Q
                           => sec_df2_inst_arx_z1_reg_4_port);
   sec_df2_inst_arx_z1_reg_reg_5 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p1_5_port, CK => clock, RB => resetn, Q
                           => sec_df2_inst_arx_z1_reg_5_port);
   sec_df2_inst_arx_z2_reg_reg_6 : DFFRPQ1 port map( D => 
                           sec_df2_inst_arx_z1_reg_6_port, CK => clock, RB => 
                           resetn, Q => sec_df2_inst_arx_z2_reg_6_port);
   sec_df2_inst_arx_z1_reg_reg_6 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p1_6_port, CK => clock, RB => resetn, Q
                           => sec_df2_inst_arx_z1_reg_6_port);
   sec_df2_inst_arx_z2_reg_reg_5 : DFFRPQ1 port map( D => 
                           sec_df2_inst_arx_z1_reg_5_port, CK => clock, RB => 
                           resetn, Q => sec_df2_inst_arx_z2_reg_5_port);
   sec_df2_inst_arx_z1_reg_reg_7 : DFFRPQ1 port map( D => 
                           sec_df2_inst_p1_7_port, CK => clock, RB => resetn, Q
                           => sec_df2_inst_m2_14);
   sec_df2_inst_arx_z2_reg_reg_7 : DFFRPQ1 port map( D => sec_df2_inst_m2_14, 
                           CK => clock, RB => resetn, Q => 
                           sec_df2_inst_arx_z2_reg_7_port);
   sec_df2_inst_add_139_U1_14 : ADFULD1 port map( A => sec_df2_inst_m1_15, B =>
                           sec_df2_inst_p4_7, CI => 
                           sec_df2_inst_add_139_carry_14_port, CO => 
                           sec_df2_inst_n_1064, S => sec_df2_inst_N26);
   sec_df2_inst_add_139_U1_13 : ADFULD1 port map( A => sec_df2_inst_m1_13, B =>
                           sec_df2_inst_p4_6, CI => 
                           sec_df2_inst_add_139_carry_13_port, CO => 
                           sec_df2_inst_add_139_carry_14_port, S => 
                           sec_df2_inst_N25);
   sec_df2_inst_add_139_U1_12 : ADFULD1 port map( A => sec_df2_inst_m1_12, B =>
                           sec_df2_inst_p4_5, CI => 
                           sec_df2_inst_add_139_carry_12_port, CO => 
                           sec_df2_inst_add_139_carry_13_port, S => 
                           sec_df2_inst_N24);
   sec_df2_inst_add_139_U1_11 : ADFULD1 port map( A => sec_df2_inst_m1_11, B =>
                           sec_df2_inst_p4_4, CI => 
                           sec_df2_inst_add_139_carry_11_port, CO => 
                           sec_df2_inst_add_139_carry_12_port, S => 
                           sec_df2_inst_N23);
   sec_df2_inst_add_139_U1_10 : ADFULD1 port map( A => sec_df2_inst_m1_10, B =>
                           sec_df2_inst_p4_3, CI => 
                           sec_df2_inst_add_139_carry_10_port, CO => 
                           sec_df2_inst_add_139_carry_11_port, S => 
                           sec_df2_inst_N22);
   sec_df2_inst_add_139_U1_9 : ADFULD1 port map( A => sec_df2_inst_m1_9, B => 
                           sec_df2_inst_p4_2, CI => 
                           sec_df2_inst_add_139_carry_9_port, CO => 
                           sec_df2_inst_add_139_carry_10_port, S => 
                           sec_df2_inst_N21);
   sec_df2_inst_add_139_U1_8 : ADFULD1 port map( A => sec_df2_inst_m1_8, B => 
                           sec_df2_inst_p4_1, CI => 
                           sec_df2_inst_add_139_carry_8_port, CO => 
                           sec_df2_inst_add_139_carry_9_port, S => 
                           sec_df2_inst_N20);
   sec_df2_inst_mult_133_U2 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z2_reg_7_port, B => 
                           sec_df2_inst_n70, CI => sec_df2_inst_mult_133_n2, CO
                           => sec_df2_inst_mult_133_n1, S => sec_df2_inst_m4_13
                           );
   sec_df2_inst_mult_133_U3 : ADFULD1 port map( A => sec_df2_inst_mult_133_n15,
                           B => sec_df2_inst_arx_z2_reg_6_port, CI => 
                           sec_df2_inst_mult_133_n3, CO => 
                           sec_df2_inst_mult_133_n2, S => sec_df2_inst_m4_12);
   sec_df2_inst_mult_133_U4 : ADFULD1 port map( A => sec_df2_inst_mult_133_n16,
                           B => sec_df2_inst_mult_133_n17, CI => 
                           sec_df2_inst_mult_133_n4, CO => 
                           sec_df2_inst_mult_133_n3, S => sec_df2_inst_m4_11);
   sec_df2_inst_mult_133_U5 : ADFULD1 port map( A => sec_df2_inst_mult_133_n18,
                           B => sec_df2_inst_mult_133_n19, CI => 
                           sec_df2_inst_mult_133_n5, CO => 
                           sec_df2_inst_mult_133_n4, S => sec_df2_inst_m4_10);
   sec_df2_inst_mult_133_U6 : ADFULD1 port map( A => sec_df2_inst_mult_133_n20,
                           B => sec_df2_inst_mult_133_n21, CI => 
                           sec_df2_inst_mult_133_n6, CO => 
                           sec_df2_inst_mult_133_n5, S => sec_df2_inst_m4_9);
   sec_df2_inst_mult_133_U7 : ADFULD1 port map( A => sec_df2_inst_mult_133_n22,
                           B => sec_df2_inst_mult_133_n23, CI => 
                           sec_df2_inst_mult_133_n7, CO => 
                           sec_df2_inst_mult_133_n6, S => sec_df2_inst_m4_8);
   sec_df2_inst_mult_133_U8 : ADFULD1 port map( A => sec_df2_inst_mult_133_n24,
                           B => sec_df2_inst_mult_133_n25, CI => 
                           sec_df2_inst_mult_133_n8, CO => 
                           sec_df2_inst_mult_133_n7, S => sec_df2_inst_m4_7);
   sec_df2_inst_mult_133_U9 : ADFULD1 port map( A => sec_df2_inst_mult_133_n26,
                           B => sec_df2_inst_m5_2, CI => 
                           sec_df2_inst_mult_133_n9, CO => 
                           sec_df2_inst_mult_133_n8, S => sec_df2_inst_m4_6);
   sec_df2_inst_mult_133_U10 : ADFULD1 port map( A => sec_df2_inst_m5_1, B => 
                           sec_df2_inst_n60, CI => sec_df2_inst_mult_133_n10, 
                           CO => sec_df2_inst_mult_133_n9, S => 
                           sec_df2_inst_m4_5);
   sec_df2_inst_mult_133_U11 : ADFULD1 port map( A => sec_df2_inst_m4_0, B => 
                           sec_df2_inst_n50, CI => sec_df2_inst_mult_133_n11, 
                           CO => sec_df2_inst_mult_133_n10, S => 
                           sec_df2_inst_m4_4);
   sec_df2_inst_mult_133_U12 : ADHALFDL port map( A => 
                           sec_df2_inst_mult_133_n12, B => sec_df2_inst_n40, CO
                           => sec_df2_inst_mult_133_n11, S => sec_df2_inst_m4_3
                           );
   sec_df2_inst_mult_133_U13 : ADHALFDL port map( A => 
                           sec_df2_inst_mult_133_n13, B => sec_df2_inst_n30, CO
                           => sec_df2_inst_mult_133_n12, S => sec_df2_inst_m4_2
                           );
   sec_df2_inst_mult_133_U14 : ADHALFDL port map( A => sec_df2_inst_n110, B => 
                           sec_df2_inst_n27, CO => sec_df2_inst_mult_133_n13, S
                           => sec_df2_inst_m4_1);
   sec_df2_inst_mult_133_U16 : ADFULD1 port map( A => sec_df2_inst_n50, B => 
                           sec_df2_inst_n80, CI => sec_df2_inst_n60, CO => 
                           sec_df2_inst_mult_133_n15, S => 
                           sec_df2_inst_mult_133_n16);
   sec_df2_inst_mult_133_U17 : ADFULD1 port map( A => sec_df2_inst_n40, B => 
                           sec_df2_inst_arx_z2_reg_4_port, CI => 
                           sec_df2_inst_arx_z2_reg_6_port, CO => 
                           sec_df2_inst_mult_133_n17, S => 
                           sec_df2_inst_mult_133_n18);
   sec_df2_inst_mult_133_U18 : ADFULD1 port map( A => sec_df2_inst_n30, B => 
                           sec_df2_inst_arx_z2_reg_3_port, CI => 
                           sec_df2_inst_arx_z2_reg_5_port, CO => 
                           sec_df2_inst_mult_133_n19, S => 
                           sec_df2_inst_mult_133_n20);
   sec_df2_inst_mult_133_U19 : ADFULD1 port map( A => sec_df2_inst_n27, B => 
                           sec_df2_inst_m5_2, CI => 
                           sec_df2_inst_arx_z2_reg_4_port, CO => 
                           sec_df2_inst_mult_133_n21, S => 
                           sec_df2_inst_mult_133_n22);
   sec_df2_inst_mult_133_U20 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z2_reg_7_port, B => 
                           sec_df2_inst_m5_1, CI => 
                           sec_df2_inst_arx_z2_reg_3_port, CO => 
                           sec_df2_inst_mult_133_n23, S => 
                           sec_df2_inst_mult_133_n24);
   sec_df2_inst_mult_131_U2 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_6_port, B => 
                           sec_df2_inst_m2_14, CI => sec_df2_inst_mult_131_n2, 
                           CO => sec_df2_inst_m2_13, S => sec_df2_inst_m2_12);
   sec_df2_inst_mult_131_U3 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_5_port, B => 
                           sec_df2_inst_m2_14, CI => sec_df2_inst_mult_131_n3, 
                           CO => sec_df2_inst_mult_131_n2, S => 
                           sec_df2_inst_m2_11);
   sec_df2_inst_mult_131_U4 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_4_port, B => 
                           sec_df2_inst_m2_14, CI => sec_df2_inst_mult_131_n4, 
                           CO => sec_df2_inst_mult_131_n3, S => 
                           sec_df2_inst_m2_10);
   sec_df2_inst_mult_131_U5 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_3_port, B => 
                           sec_df2_inst_m2_14, CI => sec_df2_inst_mult_131_n5, 
                           CO => sec_df2_inst_mult_131_n4, S => 
                           sec_df2_inst_m2_9);
   sec_df2_inst_mult_131_U6 : ADFULD1 port map( A => sec_df2_inst_mult_131_n13,
                           B => sec_df2_inst_arx_z1_reg_2_port, CI => 
                           sec_df2_inst_mult_131_n6, CO => 
                           sec_df2_inst_mult_131_n5, S => sec_df2_inst_m2_8);
   sec_df2_inst_mult_131_U7 : ADFULD1 port map( A => sec_df2_inst_mult_131_n14,
                           B => sec_df2_inst_mult_131_n15, CI => 
                           sec_df2_inst_mult_131_n7, CO => 
                           sec_df2_inst_mult_131_n6, S => sec_df2_inst_m2_7);
   sec_df2_inst_mult_131_U8 : ADFULD1 port map( A => sec_df2_inst_mult_131_n16,
                           B => sec_df2_inst_m3_1, CI => 
                           sec_df2_inst_mult_131_n8, CO => 
                           sec_df2_inst_mult_131_n7, S => sec_df2_inst_m2_6);
   sec_df2_inst_mult_131_U9 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_5_port, B => 
                           sec_df2_inst_arx_z1_reg_4_port, CI => 
                           sec_df2_inst_mult_131_n9, CO => 
                           sec_df2_inst_mult_131_n8, S => sec_df2_inst_m2_5);
   sec_df2_inst_mult_131_U10 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_4_port, B => 
                           sec_df2_inst_arx_z1_reg_3_port, CI => 
                           sec_df2_inst_mult_131_n10, CO => 
                           sec_df2_inst_mult_131_n9, S => sec_df2_inst_m2_4);
   sec_df2_inst_mult_131_U11 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_3_port, B => 
                           sec_df2_inst_arx_z1_reg_2_port, CI => 
                           sec_df2_inst_mult_131_n11, CO => 
                           sec_df2_inst_mult_131_n10, S => sec_df2_inst_m2_3);
   sec_df2_inst_mult_131_U12 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_2_port, B => 
                           sec_df2_inst_m3_2, CI => sec_df2_inst_mult_131_n12, 
                           CO => sec_df2_inst_mult_131_n11, S => 
                           sec_df2_inst_m2_2);
   sec_df2_inst_mult_131_U13 : ADHALFDL port map( A => sec_df2_inst_m3_2, B => 
                           sec_df2_inst_m3_1, CO => sec_df2_inst_mult_131_n12, 
                           S => sec_df2_inst_m2_1);
   sec_df2_inst_mult_131_U14 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_6_port, B => 
                           sec_df2_inst_m2_14, CI => sec_df2_inst_m3_2, CO => 
                           sec_df2_inst_mult_131_n13, S => 
                           sec_df2_inst_mult_131_n14);
   sec_df2_inst_mult_131_U15 : ADHALFDL port map( A => 
                           sec_df2_inst_arx_z1_reg_5_port, B => 
                           sec_df2_inst_arx_z1_reg_6_port, CO => 
                           sec_df2_inst_mult_131_n15, S => 
                           sec_df2_inst_mult_131_n16);
   sec_df2_inst_mult_134_U2 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z2_reg_6_port, B => 
                           sec_df2_inst_n80, CI => sec_df2_inst_mult_134_n2, CO
                           => sec_df2_inst_mult_134_n1, S => sec_df2_inst_m5_13
                           );
   sec_df2_inst_mult_134_U3 : ADFULD1 port map( A => sec_df2_inst_n70, B => 
                           sec_df2_inst_arx_z2_reg_5_port, CI => 
                           sec_df2_inst_mult_134_n3, CO => 
                           sec_df2_inst_mult_134_n2, S => sec_df2_inst_m5_12);
   sec_df2_inst_mult_134_U4 : ADFULD1 port map( A => sec_df2_inst_mult_134_n16,
                           B => sec_df2_inst_n60, CI => 
                           sec_df2_inst_mult_134_n4, CO => 
                           sec_df2_inst_mult_134_n3, S => sec_df2_inst_m5_11);
   sec_df2_inst_mult_134_U5 : ADFULD1 port map( A => sec_df2_inst_mult_134_n17,
                           B => sec_df2_inst_mult_134_n18, CI => 
                           sec_df2_inst_mult_134_n5, CO => 
                           sec_df2_inst_mult_134_n4, S => sec_df2_inst_m5_10);
   sec_df2_inst_mult_134_U6 : ADFULD1 port map( A => sec_df2_inst_mult_134_n19,
                           B => sec_df2_inst_mult_134_n20, CI => 
                           sec_df2_inst_mult_134_n6, CO => 
                           sec_df2_inst_mult_134_n5, S => sec_df2_inst_m5_9);
   sec_df2_inst_mult_134_U7 : ADFULD1 port map( A => sec_df2_inst_mult_134_n21,
                           B => sec_df2_inst_mult_134_n22, CI => 
                           sec_df2_inst_mult_134_n7, CO => 
                           sec_df2_inst_mult_134_n6, S => sec_df2_inst_m5_8);
   sec_df2_inst_mult_134_U8 : ADFULD1 port map( A => sec_df2_inst_mult_134_n23,
                           B => sec_df2_inst_mult_134_n24, CI => 
                           sec_df2_inst_mult_134_n8, CO => 
                           sec_df2_inst_mult_134_n7, S => sec_df2_inst_m5_7);
   sec_df2_inst_mult_134_U9 : ADFULD1 port map( A => sec_df2_inst_mult_134_n25,
                           B => sec_df2_inst_m4_0, CI => 
                           sec_df2_inst_mult_134_n9, CO => 
                           sec_df2_inst_mult_134_n8, S => sec_df2_inst_m5_6);
   sec_df2_inst_mult_134_U10 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z2_reg_5_port, B => 
                           sec_df2_inst_n30, CI => sec_df2_inst_mult_134_n10, 
                           CO => sec_df2_inst_mult_134_n9, S => 
                           sec_df2_inst_m5_5);
   sec_df2_inst_mult_134_U11 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z2_reg_4_port, B => 
                           sec_df2_inst_n27, CI => sec_df2_inst_mult_134_n11, 
                           CO => sec_df2_inst_mult_134_n10, S => 
                           sec_df2_inst_m5_4);
   sec_df2_inst_mult_134_U16 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z2_reg_7_port, B => 
                           sec_df2_inst_n70, CI => 
                           sec_df2_inst_arx_z2_reg_4_port, CO => 
                           sec_df2_inst_mult_134_n16, S => 
                           sec_df2_inst_mult_134_n17);
   sec_df2_inst_mult_134_U17 : ADFULD1 port map( A => sec_df2_inst_n60, B => 
                           sec_df2_inst_arx_z2_reg_6_port, CI => 
                           sec_df2_inst_arx_z2_reg_3_port, CO => 
                           sec_df2_inst_mult_134_n18, S => 
                           sec_df2_inst_mult_134_n19);
   sec_df2_inst_mult_134_U18 : ADFULD1 port map( A => sec_df2_inst_n80, B => 
                           sec_df2_inst_arx_z2_reg_5_port, CI => 
                           sec_df2_inst_m5_2, CO => sec_df2_inst_mult_134_n20, 
                           S => sec_df2_inst_mult_134_n21);
   sec_df2_inst_mult_134_U19 : ADFULD1 port map( A => sec_df2_inst_n50, B => 
                           sec_df2_inst_arx_z2_reg_7_port, CI => 
                           sec_df2_inst_m5_1, CO => sec_df2_inst_mult_134_n22, 
                           S => sec_df2_inst_mult_134_n23);
   sec_df2_inst_mult_134_U20 : ADHALFDL port map( A => 
                           sec_df2_inst_arx_z2_reg_6_port, B => 
                           sec_df2_inst_n40, CO => sec_df2_inst_mult_134_n24, S
                           => sec_df2_inst_mult_134_n25);
   sec_df2_inst_add_1_root_add_136_U1_7 : EXOR3D1 port map( A1 => 
                           sec_df2_inst_N8, A2 => data_in(7), A3 => 
                           sec_df2_inst_add_1_root_add_136_carry_7_port, Z => 
                           sec_df2_inst_p1_7_port);
   sec_df2_inst_add_1_root_add_136_U1_0 : ADFULD1 port map( A => 
                           sec_df2_inst_N1, B => data_in(0), CI => 
                           sec_df2_inst_N0, CO => 
                           sec_df2_inst_add_1_root_add_136_carry_1_port, S => 
                           sec_df2_inst_p1_0_port);
   sec_df2_inst_add_1_root_add_136_U1_1 : ADFULD1 port map( A => 
                           sec_df2_inst_N2, B => data_in(1), CI => 
                           sec_df2_inst_add_1_root_add_136_carry_1_port, CO => 
                           sec_df2_inst_add_1_root_add_136_carry_2_port, S => 
                           sec_df2_inst_p1_1_port);
   sec_df2_inst_add_1_root_add_136_U1_2 : ADFULD1 port map( A => 
                           sec_df2_inst_N3, B => data_in(2), CI => 
                           sec_df2_inst_add_1_root_add_136_carry_2_port, CO => 
                           sec_df2_inst_add_1_root_add_136_carry_3_port, S => 
                           sec_df2_inst_p1_2_port);
   sec_df2_inst_add_1_root_add_136_U1_3 : ADFULD1 port map( A => 
                           sec_df2_inst_N4, B => data_in(3), CI => 
                           sec_df2_inst_add_1_root_add_136_carry_3_port, CO => 
                           sec_df2_inst_add_1_root_add_136_carry_4_port, S => 
                           sec_df2_inst_p1_3_port);
   sec_df2_inst_add_1_root_add_136_U1_4 : ADFULD1 port map( A => 
                           sec_df2_inst_N5, B => data_in(4), CI => 
                           sec_df2_inst_add_1_root_add_136_carry_4_port, CO => 
                           sec_df2_inst_add_1_root_add_136_carry_5_port, S => 
                           sec_df2_inst_p1_4_port);
   sec_df2_inst_add_1_root_add_136_U1_5 : ADFULD1 port map( A => 
                           sec_df2_inst_N6, B => data_in(5), CI => 
                           sec_df2_inst_add_1_root_add_136_carry_5_port, CO => 
                           sec_df2_inst_add_1_root_add_136_carry_6_port, S => 
                           sec_df2_inst_p1_5_port);
   sec_df2_inst_add_1_root_add_136_U1_6 : ADFULD1 port map( A => 
                           sec_df2_inst_N7, B => data_in(6), CI => 
                           sec_df2_inst_add_1_root_add_136_carry_6_port, CO => 
                           sec_df2_inst_add_1_root_add_136_carry_7_port, S => 
                           sec_df2_inst_p1_6_port);
   sec_df2_inst_mult_137_U47 : NAN2D1 port map( A1 => sec_df2_inst_p1_0_port, 
                           A2 => sec_df2_inst_mult_137_n72, Z => 
                           sec_df2_inst_mult_137_n78);
   sec_df2_inst_mult_137_U46 : NAN2D1 port map( A1 => sec_df2_inst_mult_137_n78
                           , A2 => sec_df2_inst_p1_4_port, Z => 
                           sec_df2_inst_mult_137_n76);
   sec_df2_inst_mult_137_U45 : NAN2M1D1 port map( A1 => sec_df2_inst_p1_1_port,
                           A2 => sec_df2_inst_mult_137_n78, Z => 
                           sec_df2_inst_mult_137_n77);
   sec_df2_inst_mult_137_U44 : OAI211D1 port map( A1 => sec_df2_inst_p1_1_port,
                           A2 => sec_df2_inst_mult_137_n71, B => 
                           sec_df2_inst_mult_137_n76, C => 
                           sec_df2_inst_mult_137_n77, Z => 
                           sec_df2_inst_mult_137_n75);
   sec_df2_inst_mult_137_U43 : NAN2D1 port map( A1 => sec_df2_inst_mult_137_n75
                           , A2 => sec_df2_inst_p1_5_port, Z => 
                           sec_df2_inst_mult_137_n73);
   sec_df2_inst_mult_137_U42 : NAN2M1D1 port map( A1 => sec_df2_inst_p1_2_port,
                           A2 => sec_df2_inst_mult_137_n75, Z => 
                           sec_df2_inst_mult_137_n74);
   sec_df2_inst_mult_137_U41 : OAI211D1 port map( A1 => sec_df2_inst_p1_2_port,
                           A2 => sec_df2_inst_mult_137_n70, B => 
                           sec_df2_inst_mult_137_n73, C => 
                           sec_df2_inst_mult_137_n74, Z => 
                           sec_df2_inst_mult_137_n9);
   sec_df2_inst_mult_137_U40 : INVD1 port map( A => sec_df2_inst_p1_6_port, Z 
                           => sec_df2_inst_mult_137_n69);
   sec_df2_inst_mult_137_U39 : INVD1 port map( A => sec_df2_inst_p1_3_port, Z 
                           => sec_df2_inst_mult_137_n72);
   sec_df2_inst_mult_137_U38 : INVD1 port map( A => sec_df2_inst_p1_4_port, Z 
                           => sec_df2_inst_mult_137_n71);
   sec_df2_inst_mult_137_U37 : INVD1 port map( A => sec_df2_inst_p1_5_port, Z 
                           => sec_df2_inst_mult_137_n70);
   sec_df2_inst_mult_137_U36 : INVD1 port map( A => sec_df2_inst_p1_7_port, Z 
                           => sec_df2_inst_mult_137_n68);
   sec_df2_inst_mult_137_U35 : INVD1 port map( A => sec_df2_inst_mult_137_n1, Z
                           => sec_df2_inst_m1_15);
   sec_df2_inst_mult_137_U20 : ADHALFDL port map( A => sec_df2_inst_p1_6_port, 
                           B => sec_df2_inst_mult_137_n72, CO => 
                           sec_df2_inst_mult_137_n24, S => 
                           sec_df2_inst_mult_137_n25);
   sec_df2_inst_mult_137_U19 : ADFULD1 port map( A => sec_df2_inst_mult_137_n71
                           , B => sec_df2_inst_p1_7_port, CI => 
                           sec_df2_inst_p1_1_port, CO => 
                           sec_df2_inst_mult_137_n22, S => 
                           sec_df2_inst_mult_137_n23);
   sec_df2_inst_mult_137_U18 : ADFULD1 port map( A => sec_df2_inst_mult_137_n68
                           , B => sec_df2_inst_p1_5_port, CI => 
                           sec_df2_inst_p1_2_port, CO => 
                           sec_df2_inst_mult_137_n20, S => 
                           sec_df2_inst_mult_137_n21);
   sec_df2_inst_mult_137_U17 : ADFULD1 port map( A => sec_df2_inst_mult_137_n70
                           , B => sec_df2_inst_p1_6_port, CI => 
                           sec_df2_inst_p1_3_port, CO => 
                           sec_df2_inst_mult_137_n18, S => 
                           sec_df2_inst_mult_137_n19);
   sec_df2_inst_mult_137_U16 : ADFULD1 port map( A => sec_df2_inst_p1_7_port, B
                           => sec_df2_inst_mult_137_n69, CI => 
                           sec_df2_inst_p1_4_port, CO => 
                           sec_df2_inst_mult_137_n16, S => 
                           sec_df2_inst_mult_137_n17);
   sec_df2_inst_mult_137_U9 : ADFULD1 port map( A => sec_df2_inst_mult_137_n25,
                           B => sec_df2_inst_p1_0_port, CI => 
                           sec_df2_inst_mult_137_n9, CO => 
                           sec_df2_inst_mult_137_n8, S => sec_df2_inst_N18);
   sec_df2_inst_mult_137_U8 : ADFULD1 port map( A => sec_df2_inst_mult_137_n23,
                           B => sec_df2_inst_mult_137_n24, CI => 
                           sec_df2_inst_mult_137_n8, CO => 
                           sec_df2_inst_mult_137_n7, S => sec_df2_inst_m1_7);
   sec_df2_inst_mult_137_U7 : ADFULD1 port map( A => sec_df2_inst_mult_137_n21,
                           B => sec_df2_inst_mult_137_n22, CI => 
                           sec_df2_inst_mult_137_n7, CO => 
                           sec_df2_inst_mult_137_n6, S => sec_df2_inst_m1_8);
   sec_df2_inst_mult_137_U6 : ADFULD1 port map( A => sec_df2_inst_mult_137_n19,
                           B => sec_df2_inst_mult_137_n20, CI => 
                           sec_df2_inst_mult_137_n6, CO => 
                           sec_df2_inst_mult_137_n5, S => sec_df2_inst_m1_9);
   sec_df2_inst_mult_137_U5 : ADFULD1 port map( A => sec_df2_inst_mult_137_n17,
                           B => sec_df2_inst_mult_137_n18, CI => 
                           sec_df2_inst_mult_137_n5, CO => 
                           sec_df2_inst_mult_137_n4, S => sec_df2_inst_m1_10);
   sec_df2_inst_mult_137_U4 : ADFULD1 port map( A => sec_df2_inst_mult_137_n16,
                           B => sec_df2_inst_mult_137_n70, CI => 
                           sec_df2_inst_mult_137_n4, CO => 
                           sec_df2_inst_mult_137_n3, S => sec_df2_inst_m1_11);
   sec_df2_inst_mult_137_U3 : ADFULD1 port map( A => sec_df2_inst_mult_137_n69,
                           B => sec_df2_inst_p1_5_port, CI => 
                           sec_df2_inst_mult_137_n3, CO => 
                           sec_df2_inst_mult_137_n2, S => sec_df2_inst_m1_12);
   sec_df2_inst_mult_137_U2 : ADFULD1 port map( A => sec_df2_inst_p1_6_port, B 
                           => sec_df2_inst_mult_137_n68, CI => 
                           sec_df2_inst_mult_137_n2, CO => 
                           sec_df2_inst_mult_137_n1, S => sec_df2_inst_m1_13);
   sec_df2_inst_add_135_U10 : OAI211D1 port map( A1 => sec_df2_inst_m2_1, A2 =>
                           sec_df2_inst_m4_1, B => sec_df2_inst_m3_1, C => 
                           sec_df2_inst_m4_0, Z => sec_df2_inst_add_135_n9);
   sec_df2_inst_add_135_U9 : OAI21M20D1 port map( A1 => sec_df2_inst_m2_1, A2 
                           => sec_df2_inst_m4_1, B => sec_df2_inst_add_135_n9, 
                           Z => sec_df2_inst_add_135_n7);
   sec_df2_inst_add_135_U8 : OAI21D1 port map( A1 => sec_df2_inst_m2_2, A2 => 
                           sec_df2_inst_add_135_n7, B => sec_df2_inst_m4_2, Z 
                           => sec_df2_inst_add_135_n8);
   sec_df2_inst_add_135_U7 : OAI21M20D1 port map( A1 => sec_df2_inst_add_135_n7
                           , A2 => sec_df2_inst_m2_2, B => 
                           sec_df2_inst_add_135_n8, Z => 
                           sec_df2_inst_add_135_n5);
   sec_df2_inst_add_135_U6 : OAI21D1 port map( A1 => sec_df2_inst_m2_3, A2 => 
                           sec_df2_inst_add_135_n5, B => sec_df2_inst_m4_3, Z 
                           => sec_df2_inst_add_135_n6);
   sec_df2_inst_add_135_U5 : OAI21M20D1 port map( A1 => sec_df2_inst_add_135_n5
                           , A2 => sec_df2_inst_m2_3, B => 
                           sec_df2_inst_add_135_n6, Z => 
                           sec_df2_inst_add_135_n3);
   sec_df2_inst_add_135_U4 : OAI21D1 port map( A1 => sec_df2_inst_m2_4, A2 => 
                           sec_df2_inst_add_135_n3, B => sec_df2_inst_m4_4, Z 
                           => sec_df2_inst_add_135_n4);
   sec_df2_inst_add_135_U3 : OAI21M20D1 port map( A1 => sec_df2_inst_add_135_n3
                           , A2 => sec_df2_inst_m2_4, B => 
                           sec_df2_inst_add_135_n4, Z => 
                           sec_df2_inst_add_135_n1);
   sec_df2_inst_add_135_U2 : OAI21D1 port map( A1 => sec_df2_inst_m2_5, A2 => 
                           sec_df2_inst_add_135_n1, B => sec_df2_inst_m4_5, Z 
                           => sec_df2_inst_add_135_n2);
   sec_df2_inst_add_135_U1 : OAI21M20D1 port map( A1 => sec_df2_inst_add_135_n1
                           , A2 => sec_df2_inst_m2_5, B => 
                           sec_df2_inst_add_135_n2, Z => 
                           sec_df2_inst_add_135_carry_6_port);
   sec_df2_inst_add_135_U1_14 : EXOR3D1 port map( A1 => sec_df2_inst_m2_14, A2 
                           => sec_df2_inst_m4_15, A3 => 
                           sec_df2_inst_add_135_carry_14_port, Z => 
                           sec_df2_inst_N8);
   sec_df2_inst_add_135_U1_6 : ADFULD1 port map( A => sec_df2_inst_m2_6, B => 
                           sec_df2_inst_m4_6, CI => 
                           sec_df2_inst_add_135_carry_6_port, CO => 
                           sec_df2_inst_add_135_carry_7_port, S => 
                           sec_df2_inst_N0);
   sec_df2_inst_add_135_U1_7 : ADFULD1 port map( A => sec_df2_inst_m2_7, B => 
                           sec_df2_inst_m4_7, CI => 
                           sec_df2_inst_add_135_carry_7_port, CO => 
                           sec_df2_inst_add_135_carry_8_port, S => 
                           sec_df2_inst_N1);
   sec_df2_inst_add_135_U1_8 : ADFULD1 port map( A => sec_df2_inst_m2_8, B => 
                           sec_df2_inst_m4_8, CI => 
                           sec_df2_inst_add_135_carry_8_port, CO => 
                           sec_df2_inst_add_135_carry_9_port, S => 
                           sec_df2_inst_N2);
   sec_df2_inst_add_135_U1_9 : ADFULD1 port map( A => sec_df2_inst_m2_9, B => 
                           sec_df2_inst_m4_9, CI => 
                           sec_df2_inst_add_135_carry_9_port, CO => 
                           sec_df2_inst_add_135_carry_10_port, S => 
                           sec_df2_inst_N3);
   sec_df2_inst_add_135_U1_10 : ADFULD1 port map( A => sec_df2_inst_m2_10, B =>
                           sec_df2_inst_m4_10, CI => 
                           sec_df2_inst_add_135_carry_10_port, CO => 
                           sec_df2_inst_add_135_carry_11_port, S => 
                           sec_df2_inst_N4);
   sec_df2_inst_add_135_U1_11 : ADFULD1 port map( A => sec_df2_inst_m2_11, B =>
                           sec_df2_inst_m4_11, CI => 
                           sec_df2_inst_add_135_carry_11_port, CO => 
                           sec_df2_inst_add_135_carry_12_port, S => 
                           sec_df2_inst_N5);
   sec_df2_inst_add_135_U1_12 : ADFULD1 port map( A => sec_df2_inst_m2_12, B =>
                           sec_df2_inst_m4_12, CI => 
                           sec_df2_inst_add_135_carry_12_port, CO => 
                           sec_df2_inst_add_135_carry_13_port, S => 
                           sec_df2_inst_N6);
   sec_df2_inst_add_135_U1_13 : ADFULD1 port map( A => sec_df2_inst_m2_13, B =>
                           sec_df2_inst_m4_13, CI => 
                           sec_df2_inst_add_135_carry_13_port, CO => 
                           sec_df2_inst_add_135_carry_14_port, S => 
                           sec_df2_inst_N7);
   sec_df2_inst_mult_132_U51 : NAN2D1 port map( A1 => sec_df2_inst_m3_1, A2 => 
                           sec_df2_inst_mult_132_n84, Z => 
                           sec_df2_inst_mult_132_n29);
   sec_df2_inst_mult_132_U50 : EXOR2D1 port map( A1 => 
                           sec_df2_inst_arx_z1_reg_6_port, A2 => 
                           sec_df2_inst_m3_1, Z => sec_df2_inst_mult_132_n30);
   sec_df2_inst_mult_132_U49 : EXOR3D1 port map( A1 => sec_df2_inst_mult_132_n2
                           , A2 => sec_df2_inst_m2_14, A3 => 
                           sec_df2_inst_mult_132_n84, Z => sec_df2_inst_m3_14);
   sec_df2_inst_mult_132_U48 : INVD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_4_port, Z => 
                           sec_df2_inst_mult_132_n86);
   sec_df2_inst_mult_132_U47 : INVD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_2_port, Z => 
                           sec_df2_inst_mult_132_n88);
   sec_df2_inst_mult_132_U46 : INVD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_3_port, Z => 
                           sec_df2_inst_mult_132_n87);
   sec_df2_inst_mult_132_U45 : INVD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_6_port, Z => 
                           sec_df2_inst_mult_132_n84);
   sec_df2_inst_mult_132_U44 : INVD1 port map( A => sec_df2_inst_m2_14, Z => 
                           sec_df2_inst_mult_132_n83);
   sec_df2_inst_mult_132_U43 : INVD1 port map( A => sec_df2_inst_m3_2, Z => 
                           sec_df2_inst_mult_132_n89);
   sec_df2_inst_mult_132_U42 : INVD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_5_port, Z => 
                           sec_df2_inst_mult_132_n85);
   sec_df2_inst_mult_132_U26 : ADHALFDL port map( A => sec_df2_inst_m3_2, B => 
                           sec_df2_inst_arx_z1_reg_3_port, CO => 
                           sec_df2_inst_mult_132_n35, S => 
                           sec_df2_inst_mult_132_n36);
   sec_df2_inst_mult_132_U25 : ADFULD1 port map( A => sec_df2_inst_m3_2, B => 
                           sec_df2_inst_arx_z1_reg_4_port, CI => 
                           sec_df2_inst_arx_z1_reg_2_port, CO => 
                           sec_df2_inst_mult_132_n33, S => 
                           sec_df2_inst_mult_132_n34);
   sec_df2_inst_mult_132_U24 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_2_port, B => 
                           sec_df2_inst_arx_z1_reg_5_port, CI => 
                           sec_df2_inst_arx_z1_reg_3_port, CO => 
                           sec_df2_inst_mult_132_n31, S => 
                           sec_df2_inst_mult_132_n32);
   sec_df2_inst_mult_132_U21 : ADFULD1 port map( A => 
                           sec_df2_inst_arx_z1_reg_3_port, B => 
                           sec_df2_inst_arx_z1_reg_4_port, CI => 
                           sec_df2_inst_mult_132_n30, CO => 
                           sec_df2_inst_mult_132_n27, S => 
                           sec_df2_inst_mult_132_n28);
   sec_df2_inst_mult_132_U20 : ADFULD1 port map( A => sec_df2_inst_mult_132_n89
                           , B => sec_df2_inst_m2_14, CI => 
                           sec_df2_inst_arx_z1_reg_5_port, CO => 
                           sec_df2_inst_mult_132_n25, S => 
                           sec_df2_inst_mult_132_n26);
   sec_df2_inst_mult_132_U19 : ADFULD1 port map( A => sec_df2_inst_mult_132_n29
                           , B => sec_df2_inst_arx_z1_reg_4_port, CI => 
                           sec_df2_inst_mult_132_n26, CO => 
                           sec_df2_inst_mult_132_n23, S => 
                           sec_df2_inst_mult_132_n24);
   sec_df2_inst_mult_132_U18 : ADFULD1 port map( A => sec_df2_inst_mult_132_n83
                           , B => sec_df2_inst_arx_z1_reg_2_port, CI => 
                           sec_df2_inst_arx_z1_reg_6_port, CO => 
                           sec_df2_inst_mult_132_n21, S => 
                           sec_df2_inst_mult_132_n22);
   sec_df2_inst_mult_132_U17 : ADFULD1 port map( A => sec_df2_inst_mult_132_n25
                           , B => sec_df2_inst_arx_z1_reg_5_port, CI => 
                           sec_df2_inst_mult_132_n22, CO => 
                           sec_df2_inst_mult_132_n19, S => 
                           sec_df2_inst_mult_132_n20);
   sec_df2_inst_mult_132_U16 : ADFULD1 port map( A => sec_df2_inst_mult_132_n88
                           , B => sec_df2_inst_mult_132_n87, CI => 
                           sec_df2_inst_arx_z1_reg_6_port, CO => 
                           sec_df2_inst_mult_132_n17, S => 
                           sec_df2_inst_mult_132_n18);
   sec_df2_inst_mult_132_U15 : ADFULD1 port map( A => sec_df2_inst_mult_132_n21
                           , B => sec_df2_inst_mult_132_n83, CI => 
                           sec_df2_inst_mult_132_n18, CO => 
                           sec_df2_inst_mult_132_n15, S => 
                           sec_df2_inst_mult_132_n16);
   sec_df2_inst_mult_132_U14 : ADFULD1 port map( A => sec_df2_inst_mult_132_n86
                           , B => sec_df2_inst_mult_132_n83, CI => 
                           sec_df2_inst_mult_132_n17, CO => 
                           sec_df2_inst_mult_132_n13, S => 
                           sec_df2_inst_mult_132_n14);
   sec_df2_inst_mult_132_U13 : ADHALFDL port map( A => 
                           sec_df2_inst_arx_z1_reg_2_port, B => 
                           sec_df2_inst_m3_1, CO => sec_df2_inst_mult_132_n12, 
                           S => sec_df2_inst_m3_3);
   sec_df2_inst_mult_132_U12 : ADFULD1 port map( A => sec_df2_inst_mult_132_n12
                           , B => sec_df2_inst_m3_1, CI => 
                           sec_df2_inst_mult_132_n36, CO => 
                           sec_df2_inst_mult_132_n11, S => sec_df2_inst_m3_4);
   sec_df2_inst_mult_132_U11 : ADFULD1 port map( A => sec_df2_inst_mult_132_n34
                           , B => sec_df2_inst_mult_132_n35, CI => 
                           sec_df2_inst_mult_132_n11, CO => 
                           sec_df2_inst_mult_132_n10, S => sec_df2_inst_m3_5);
   sec_df2_inst_mult_132_U10 : ADFULD1 port map( A => sec_df2_inst_mult_132_n32
                           , B => sec_df2_inst_mult_132_n33, CI => 
                           sec_df2_inst_mult_132_n10, CO => 
                           sec_df2_inst_mult_132_n9, S => sec_df2_inst_m3_6);
   sec_df2_inst_mult_132_U9 : ADFULD1 port map( A => sec_df2_inst_mult_132_n28,
                           B => sec_df2_inst_mult_132_n31, CI => 
                           sec_df2_inst_mult_132_n9, CO => 
                           sec_df2_inst_mult_132_n8, S => sec_df2_inst_m3_7);
   sec_df2_inst_mult_132_U8 : ADFULD1 port map( A => sec_df2_inst_mult_132_n24,
                           B => sec_df2_inst_mult_132_n27, CI => 
                           sec_df2_inst_mult_132_n8, CO => 
                           sec_df2_inst_mult_132_n7, S => sec_df2_inst_m3_8);
   sec_df2_inst_mult_132_U7 : ADFULD1 port map( A => sec_df2_inst_mult_132_n20,
                           B => sec_df2_inst_mult_132_n23, CI => 
                           sec_df2_inst_mult_132_n7, CO => 
                           sec_df2_inst_mult_132_n6, S => sec_df2_inst_m3_9);
   sec_df2_inst_mult_132_U6 : ADFULD1 port map( A => sec_df2_inst_mult_132_n16,
                           B => sec_df2_inst_mult_132_n19, CI => 
                           sec_df2_inst_mult_132_n6, CO => 
                           sec_df2_inst_mult_132_n5, S => sec_df2_inst_m3_10);
   sec_df2_inst_mult_132_U5 : ADFULD1 port map( A => sec_df2_inst_mult_132_n14,
                           B => sec_df2_inst_mult_132_n15, CI => 
                           sec_df2_inst_mult_132_n5, CO => 
                           sec_df2_inst_mult_132_n4, S => sec_df2_inst_m3_11);
   sec_df2_inst_mult_132_U4 : ADFULD1 port map( A => sec_df2_inst_mult_132_n13,
                           B => sec_df2_inst_arx_z1_reg_5_port, CI => 
                           sec_df2_inst_mult_132_n4, CO => 
                           sec_df2_inst_mult_132_n3, S => sec_df2_inst_m3_12);
   sec_df2_inst_mult_132_U3 : ADFULD1 port map( A => sec_df2_inst_mult_132_n85,
                           B => sec_df2_inst_arx_z1_reg_6_port, CI => 
                           sec_df2_inst_mult_132_n3, CO => 
                           sec_df2_inst_mult_132_n2, S => sec_df2_inst_m3_13);
   sec_df2_inst_add_138_U9 : OAI21D1 port map( A1 => sec_df2_inst_m3_2, A2 => 
                           sec_df2_inst_add_138_n7, B => sec_df2_inst_m5_2, Z 
                           => sec_df2_inst_add_138_n8);
   sec_df2_inst_add_138_U8 : OAI21M20D1 port map( A1 => sec_df2_inst_add_138_n7
                           , A2 => sec_df2_inst_m3_2, B => 
                           sec_df2_inst_add_138_n8, Z => 
                           sec_df2_inst_add_138_n5);
   sec_df2_inst_add_138_U7 : OAI21D1 port map( A1 => sec_df2_inst_m3_3, A2 => 
                           sec_df2_inst_add_138_n5, B => sec_df2_inst_m5_3, Z 
                           => sec_df2_inst_add_138_n6);
   sec_df2_inst_add_138_U6 : OAI21M20D1 port map( A1 => sec_df2_inst_add_138_n5
                           , A2 => sec_df2_inst_m3_3, B => 
                           sec_df2_inst_add_138_n6, Z => 
                           sec_df2_inst_add_138_n3);
   sec_df2_inst_add_138_U5 : OAI21D1 port map( A1 => sec_df2_inst_m3_4, A2 => 
                           sec_df2_inst_add_138_n3, B => sec_df2_inst_m5_4, Z 
                           => sec_df2_inst_add_138_n4);
   sec_df2_inst_add_138_U4 : OAI21M20D1 port map( A1 => sec_df2_inst_add_138_n3
                           , A2 => sec_df2_inst_m3_4, B => 
                           sec_df2_inst_add_138_n4, Z => 
                           sec_df2_inst_add_138_n1);
   sec_df2_inst_add_138_U3 : OAI21D1 port map( A1 => sec_df2_inst_m3_5, A2 => 
                           sec_df2_inst_add_138_n1, B => sec_df2_inst_m5_5, Z 
                           => sec_df2_inst_add_138_n2);
   sec_df2_inst_add_138_U2 : OAI21M20D1 port map( A1 => sec_df2_inst_add_138_n1
                           , A2 => sec_df2_inst_m3_5, B => 
                           sec_df2_inst_add_138_n2, Z => 
                           sec_df2_inst_add_138_carry_6_port);
   sec_df2_inst_add_138_U1 : AND2D1 port map( A1 => sec_df2_inst_m3_1, A2 => 
                           sec_df2_inst_m5_1, Z => sec_df2_inst_add_138_n7);
   sec_df2_inst_add_138_U1_14 : EXOR3D1 port map( A1 => sec_df2_inst_m3_14, A2 
                           => sec_df2_inst_m5_15, A3 => 
                           sec_df2_inst_add_138_carry_14_port, Z => 
                           sec_df2_inst_N17);
   sec_df2_inst_add_138_U1_6 : ADFULD1 port map( A => sec_df2_inst_m3_6, B => 
                           sec_df2_inst_m5_6, CI => 
                           sec_df2_inst_add_138_carry_6_port, CO => 
                           sec_df2_inst_add_138_carry_7_port, S => 
                           sec_df2_inst_N9);
   sec_df2_inst_add_138_U1_7 : ADFULD1 port map( A => sec_df2_inst_m3_7, B => 
                           sec_df2_inst_m5_7, CI => 
                           sec_df2_inst_add_138_carry_7_port, CO => 
                           sec_df2_inst_add_138_carry_8_port, S => 
                           sec_df2_inst_N10);
   sec_df2_inst_add_138_U1_8 : ADFULD1 port map( A => sec_df2_inst_m3_8, B => 
                           sec_df2_inst_m5_8, CI => 
                           sec_df2_inst_add_138_carry_8_port, CO => 
                           sec_df2_inst_add_138_carry_9_port, S => 
                           sec_df2_inst_N11);
   sec_df2_inst_add_138_U1_9 : ADFULD1 port map( A => sec_df2_inst_m3_9, B => 
                           sec_df2_inst_m5_9, CI => 
                           sec_df2_inst_add_138_carry_9_port, CO => 
                           sec_df2_inst_add_138_carry_10_port, S => 
                           sec_df2_inst_N12);
   sec_df2_inst_add_138_U1_10 : ADFULD1 port map( A => sec_df2_inst_m3_10, B =>
                           sec_df2_inst_m5_10, CI => 
                           sec_df2_inst_add_138_carry_10_port, CO => 
                           sec_df2_inst_add_138_carry_11_port, S => 
                           sec_df2_inst_N13);
   sec_df2_inst_add_138_U1_11 : ADFULD1 port map( A => sec_df2_inst_m3_11, B =>
                           sec_df2_inst_m5_11, CI => 
                           sec_df2_inst_add_138_carry_11_port, CO => 
                           sec_df2_inst_add_138_carry_12_port, S => 
                           sec_df2_inst_N14);
   sec_df2_inst_add_138_U1_12 : ADFULD1 port map( A => sec_df2_inst_m3_12, B =>
                           sec_df2_inst_m5_12, CI => 
                           sec_df2_inst_add_138_carry_12_port, CO => 
                           sec_df2_inst_add_138_carry_13_port, S => 
                           sec_df2_inst_N15);
   sec_df2_inst_add_138_U1_13 : ADFULD1 port map( A => sec_df2_inst_m3_13, B =>
                           sec_df2_inst_m5_13, CI => 
                           sec_df2_inst_add_138_carry_13_port, CO => 
                           sec_df2_inst_add_138_carry_14_port, S => 
                           sec_df2_inst_N16);

end flat_rtl_none_10;
